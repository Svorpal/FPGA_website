module neighboring_boids_LUT (
input [26:0] neighboring_boids,
output signed [26:0] neighboring_boids_val_out
);

reg signed [26:0] neighboring_boids_val;
assign neighboring_boids_val_out = neighboring_boids_val ;
always@(neighboring_boids) begin
    case(neighboring_boids)
        27'b000000000001000000000000000: neighboring_boids_val = 27'b000000000001000000000000000 ; // (1/1) or 1.00000000
        27'b000000000010000000000000000: neighboring_boids_val = 27'b000000000000100000000000000 ; // (1/2) or 0.50000000
        27'b000000000011000000000000000: neighboring_boids_val = 27'b000000000000010101010101010 ; // (1/3) or 0.33333333
        27'b000000000100000000000000000: neighboring_boids_val = 27'b000000000000010000000000000 ; // (1/4) or 0.25000000
        27'b000000000101000000000000000: neighboring_boids_val = 27'b000000000000001100110011001 ; // (1/5) or 0.20000000
        27'b000000000110000000000000000: neighboring_boids_val = 27'b000000000000001010101010101 ; // (1/6) or 0.16666667
        27'b000000000111000000000000000: neighboring_boids_val = 27'b000000000000001001001001001 ; // (1/7) or 0.14285714
        27'b000000001000000000000000000: neighboring_boids_val = 27'b000000000000001000000000000 ; // (1/8) or 0.12500000
        27'b000000001001000000000000000: neighboring_boids_val = 27'b000000000000000111000111000 ; // (1/9) or 0.11111111
        27'b000000001010000000000000000: neighboring_boids_val = 27'b000000000000000110011001100 ; // (1/10) or 0.10000000
        27'b000000001011000000000000000: neighboring_boids_val = 27'b000000000000000101110100010 ; // (1/11) or 0.09090909
        27'b000000001100000000000000000: neighboring_boids_val = 27'b000000000000000101010101010 ; // (1/12) or 0.08333333
        27'b000000001101000000000000000: neighboring_boids_val = 27'b000000000000000100111011000 ; // (1/13) or 0.07692308
        27'b000000001110000000000000000: neighboring_boids_val = 27'b000000000000000100100100100 ; // (1/14) or 0.07142857
        27'b000000001111000000000000000: neighboring_boids_val = 27'b000000000000000100010001000 ; // (1/15) or 0.06666667
        27'b000000010000000000000000000: neighboring_boids_val = 27'b000000000000000100000000000 ; // (1/16) or 0.06250000
        27'b000000010001000000000000000: neighboring_boids_val = 27'b000000000000000011110000111 ; // (1/17) or 0.05882353
        27'b000000010010000000000000000: neighboring_boids_val = 27'b000000000000000011100011100 ; // (1/18) or 0.05555556
        27'b000000010011000000000000000: neighboring_boids_val = 27'b000000000000000011010111100 ; // (1/19) or 0.05263158
        27'b000000010100000000000000000: neighboring_boids_val = 27'b000000000000000011001100110 ; // (1/20) or 0.05000000
        27'b000000010101000000000000000: neighboring_boids_val = 27'b000000000000000011000011000 ; // (1/21) or 0.04761905
        27'b000000010110000000000000000: neighboring_boids_val = 27'b000000000000000010111010001 ; // (1/22) or 0.04545455
        27'b000000010111000000000000000: neighboring_boids_val = 27'b000000000000000010110010000 ; // (1/23) or 0.04347826
        27'b000000011000000000000000000: neighboring_boids_val = 27'b000000000000000010101010101 ; // (1/24) or 0.04166667
        27'b000000011001000000000000000: neighboring_boids_val = 27'b000000000000000010100011110 ; // (1/25) or 0.04000000
        27'b000000011010000000000000000: neighboring_boids_val = 27'b000000000000000010011101100 ; // (1/26) or 0.03846154
        27'b000000011011000000000000000: neighboring_boids_val = 27'b000000000000000010010111101 ; // (1/27) or 0.03703704
        27'b000000011100000000000000000: neighboring_boids_val = 27'b000000000000000010010010010 ; // (1/28) or 0.03571429
        27'b000000011101000000000000000: neighboring_boids_val = 27'b000000000000000010001101001 ; // (1/29) or 0.03448276
        27'b000000011110000000000000000: neighboring_boids_val = 27'b000000000000000010001000100 ; // (1/30) or 0.03333333
        27'b000000011111000000000000000: neighboring_boids_val = 27'b000000000000000010000100001 ; // (1/31) or 0.03225806
        27'b000000100000000000000000000: neighboring_boids_val = 27'b000000000000000010000000000 ; // (1/32) or 0.03125000
        27'b000000100001000000000000000: neighboring_boids_val = 27'b000000000000000001111100000 ; // (1/33) or 0.03030303
        27'b000000100010000000000000000: neighboring_boids_val = 27'b000000000000000001111000011 ; // (1/34) or 0.02941176
        27'b000000100011000000000000000: neighboring_boids_val = 27'b000000000000000001110101000 ; // (1/35) or 0.02857143
        27'b000000100100000000000000000: neighboring_boids_val = 27'b000000000000000001110001110 ; // (1/36) or 0.02777778
        27'b000000100101000000000000000: neighboring_boids_val = 27'b000000000000000001101110101 ; // (1/37) or 0.02702703
        27'b000000100110000000000000000: neighboring_boids_val = 27'b000000000000000001101011110 ; // (1/38) or 0.02631579
        27'b000000100111000000000000000: neighboring_boids_val = 27'b000000000000000001101001000 ; // (1/39) or 0.02564103
        27'b000000101000000000000000000: neighboring_boids_val = 27'b000000000000000001100110011 ; // (1/40) or 0.02500000
        27'b000000101001000000000000000: neighboring_boids_val = 27'b000000000000000001100011111 ; // (1/41) or 0.02439024
        27'b000000101010000000000000000: neighboring_boids_val = 27'b000000000000000001100001100 ; // (1/42) or 0.02380952
        27'b000000101011000000000000000: neighboring_boids_val = 27'b000000000000000001011111010 ; // (1/43) or 0.02325581
        27'b000000101100000000000000000: neighboring_boids_val = 27'b000000000000000001011101000 ; // (1/44) or 0.02272727
        27'b000000101101000000000000000: neighboring_boids_val = 27'b000000000000000001011011000 ; // (1/45) or 0.02222222
        27'b000000101110000000000000000: neighboring_boids_val = 27'b000000000000000001011001000 ; // (1/46) or 0.02173913
        27'b000000101111000000000000000: neighboring_boids_val = 27'b000000000000000001010111001 ; // (1/47) or 0.02127660
        27'b000000110000000000000000000: neighboring_boids_val = 27'b000000000000000001010101010 ; // (1/48) or 0.02083333
        27'b000000110001000000000000000: neighboring_boids_val = 27'b000000000000000001010011100 ; // (1/49) or 0.02040816
        27'b000000110010000000000000000: neighboring_boids_val = 27'b000000000000000001010001111 ; // (1/50) or 0.02000000
        27'b000000110011000000000000000: neighboring_boids_val = 27'b000000000000000001010000010 ; // (1/51) or 0.01960784
        27'b000000110100000000000000000: neighboring_boids_val = 27'b000000000000000001001110110 ; // (1/52) or 0.01923077
        27'b000000110101000000000000000: neighboring_boids_val = 27'b000000000000000001001101010 ; // (1/53) or 0.01886792
        27'b000000110110000000000000000: neighboring_boids_val = 27'b000000000000000001001011110 ; // (1/54) or 0.01851852
        27'b000000110111000000000000000: neighboring_boids_val = 27'b000000000000000001001010011 ; // (1/55) or 0.01818182
        27'b000000111000000000000000000: neighboring_boids_val = 27'b000000000000000001001001001 ; // (1/56) or 0.01785714
        27'b000000111001000000000000000: neighboring_boids_val = 27'b000000000000000001000111110 ; // (1/57) or 0.01754386
        27'b000000111010000000000000000: neighboring_boids_val = 27'b000000000000000001000110100 ; // (1/58) or 0.01724138
        27'b000000111011000000000000000: neighboring_boids_val = 27'b000000000000000001000101011 ; // (1/59) or 0.01694915
        27'b000000111100000000000000000: neighboring_boids_val = 27'b000000000000000001000100010 ; // (1/60) or 0.01666667
        27'b000000111101000000000000000: neighboring_boids_val = 27'b000000000000000001000011001 ; // (1/61) or 0.01639344
        27'b000000111110000000000000000: neighboring_boids_val = 27'b000000000000000001000010000 ; // (1/62) or 0.01612903
        27'b000000111111000000000000000: neighboring_boids_val = 27'b000000000000000001000001000 ; // (1/63) or 0.01587302
        27'b000001000000000000000000000: neighboring_boids_val = 27'b000000000000000001000000000 ; // (1/64) or 0.01562500
        27'b000001000001000000000000000: neighboring_boids_val = 27'b000000000000000000111111000 ; // (1/65) or 0.01538462
        27'b000001000010000000000000000: neighboring_boids_val = 27'b000000000000000000111110000 ; // (1/66) or 0.01515152
        27'b000001000011000000000000000: neighboring_boids_val = 27'b000000000000000000111101001 ; // (1/67) or 0.01492537
        27'b000001000100000000000000000: neighboring_boids_val = 27'b000000000000000000111100001 ; // (1/68) or 0.01470588
        27'b000001000101000000000000000: neighboring_boids_val = 27'b000000000000000000111011010 ; // (1/69) or 0.01449275
        27'b000001000110000000000000000: neighboring_boids_val = 27'b000000000000000000111010100 ; // (1/70) or 0.01428571
        27'b000001000111000000000000000: neighboring_boids_val = 27'b000000000000000000111001101 ; // (1/71) or 0.01408451
        27'b000001001000000000000000000: neighboring_boids_val = 27'b000000000000000000111000111 ; // (1/72) or 0.01388889
        27'b000001001001000000000000000: neighboring_boids_val = 27'b000000000000000000111000000 ; // (1/73) or 0.01369863
        27'b000001001010000000000000000: neighboring_boids_val = 27'b000000000000000000110111010 ; // (1/74) or 0.01351351
        27'b000001001011000000000000000: neighboring_boids_val = 27'b000000000000000000110110100 ; // (1/75) or 0.01333333
        27'b000001001100000000000000000: neighboring_boids_val = 27'b000000000000000000110101111 ; // (1/76) or 0.01315789
        27'b000001001101000000000000000: neighboring_boids_val = 27'b000000000000000000110101001 ; // (1/77) or 0.01298701
        27'b000001001110000000000000000: neighboring_boids_val = 27'b000000000000000000110100100 ; // (1/78) or 0.01282051
        27'b000001001111000000000000000: neighboring_boids_val = 27'b000000000000000000110011110 ; // (1/79) or 0.01265823
        27'b000001010000000000000000000: neighboring_boids_val = 27'b000000000000000000110011001 ; // (1/80) or 0.01250000
        27'b000001010001000000000000000: neighboring_boids_val = 27'b000000000000000000110010100 ; // (1/81) or 0.01234568
        27'b000001010010000000000000000: neighboring_boids_val = 27'b000000000000000000110001111 ; // (1/82) or 0.01219512
        27'b000001010011000000000000000: neighboring_boids_val = 27'b000000000000000000110001010 ; // (1/83) or 0.01204819
        27'b000001010100000000000000000: neighboring_boids_val = 27'b000000000000000000110000110 ; // (1/84) or 0.01190476
        27'b000001010101000000000000000: neighboring_boids_val = 27'b000000000000000000110000001 ; // (1/85) or 0.01176471
        27'b000001010110000000000000000: neighboring_boids_val = 27'b000000000000000000101111101 ; // (1/86) or 0.01162791
        27'b000001010111000000000000000: neighboring_boids_val = 27'b000000000000000000101111000 ; // (1/87) or 0.01149425
        27'b000001011000000000000000000: neighboring_boids_val = 27'b000000000000000000101110100 ; // (1/88) or 0.01136364
        27'b000001011001000000000000000: neighboring_boids_val = 27'b000000000000000000101110000 ; // (1/89) or 0.01123596
        27'b000001011010000000000000000: neighboring_boids_val = 27'b000000000000000000101101100 ; // (1/90) or 0.01111111
        27'b000001011011000000000000000: neighboring_boids_val = 27'b000000000000000000101101000 ; // (1/91) or 0.01098901
        27'b000001011100000000000000000: neighboring_boids_val = 27'b000000000000000000101100100 ; // (1/92) or 0.01086957
        27'b000001011101000000000000000: neighboring_boids_val = 27'b000000000000000000101100000 ; // (1/93) or 0.01075269
        27'b000001011110000000000000000: neighboring_boids_val = 27'b000000000000000000101011100 ; // (1/94) or 0.01063830
        27'b000001011111000000000000000: neighboring_boids_val = 27'b000000000000000000101011000 ; // (1/95) or 0.01052632
        27'b000001100000000000000000000: neighboring_boids_val = 27'b000000000000000000101010101 ; // (1/96) or 0.01041667
        27'b000001100001000000000000000: neighboring_boids_val = 27'b000000000000000000101010001 ; // (1/97) or 0.01030928
        27'b000001100010000000000000000: neighboring_boids_val = 27'b000000000000000000101001110 ; // (1/98) or 0.01020408
        27'b000001100011000000000000000: neighboring_boids_val = 27'b000000000000000000101001010 ; // (1/99) or 0.01010101
        27'b000001100100000000000000000: neighboring_boids_val = 27'b000000000000000000101000111 ; // (1/100) or 0.01000000
        27'b000001100101000000000000000: neighboring_boids_val = 27'b000000000000000000101000100 ; // (1/101) or 0.00990099
        27'b000001100110000000000000000: neighboring_boids_val = 27'b000000000000000000101000001 ; // (1/102) or 0.00980392
        27'b000001100111000000000000000: neighboring_boids_val = 27'b000000000000000000100111110 ; // (1/103) or 0.00970874
        27'b000001101000000000000000000: neighboring_boids_val = 27'b000000000000000000100111011 ; // (1/104) or 0.00961538
        27'b000001101001000000000000000: neighboring_boids_val = 27'b000000000000000000100111000 ; // (1/105) or 0.00952381
        27'b000001101010000000000000000: neighboring_boids_val = 27'b000000000000000000100110101 ; // (1/106) or 0.00943396
        27'b000001101011000000000000000: neighboring_boids_val = 27'b000000000000000000100110010 ; // (1/107) or 0.00934579
        27'b000001101100000000000000000: neighboring_boids_val = 27'b000000000000000000100101111 ; // (1/108) or 0.00925926
        27'b000001101101000000000000000: neighboring_boids_val = 27'b000000000000000000100101100 ; // (1/109) or 0.00917431
        27'b000001101110000000000000000: neighboring_boids_val = 27'b000000000000000000100101001 ; // (1/110) or 0.00909091
        27'b000001101111000000000000000: neighboring_boids_val = 27'b000000000000000000100100111 ; // (1/111) or 0.00900901
        27'b000001110000000000000000000: neighboring_boids_val = 27'b000000000000000000100100100 ; // (1/112) or 0.00892857
        27'b000001110001000000000000000: neighboring_boids_val = 27'b000000000000000000100100001 ; // (1/113) or 0.00884956
        27'b000001110010000000000000000: neighboring_boids_val = 27'b000000000000000000100011111 ; // (1/114) or 0.00877193
        27'b000001110011000000000000000: neighboring_boids_val = 27'b000000000000000000100011100 ; // (1/115) or 0.00869565
        27'b000001110100000000000000000: neighboring_boids_val = 27'b000000000000000000100011010 ; // (1/116) or 0.00862069
        27'b000001110101000000000000000: neighboring_boids_val = 27'b000000000000000000100011000 ; // (1/117) or 0.00854701
        27'b000001110110000000000000000: neighboring_boids_val = 27'b000000000000000000100010101 ; // (1/118) or 0.00847458
        27'b000001110111000000000000000: neighboring_boids_val = 27'b000000000000000000100010011 ; // (1/119) or 0.00840336
        27'b000001111000000000000000000: neighboring_boids_val = 27'b000000000000000000100010001 ; // (1/120) or 0.00833333
        27'b000001111001000000000000000: neighboring_boids_val = 27'b000000000000000000100001110 ; // (1/121) or 0.00826446
        27'b000001111010000000000000000: neighboring_boids_val = 27'b000000000000000000100001100 ; // (1/122) or 0.00819672
        27'b000001111011000000000000000: neighboring_boids_val = 27'b000000000000000000100001010 ; // (1/123) or 0.00813008
        27'b000001111100000000000000000: neighboring_boids_val = 27'b000000000000000000100001000 ; // (1/124) or 0.00806452
        27'b000001111101000000000000000: neighboring_boids_val = 27'b000000000000000000100000110 ; // (1/125) or 0.00800000
        27'b000001111110000000000000000: neighboring_boids_val = 27'b000000000000000000100000100 ; // (1/126) or 0.00793651
        27'b000001111111000000000000000: neighboring_boids_val = 27'b000000000000000000100000010 ; // (1/127) or 0.00787402
        27'b000010000000000000000000000: neighboring_boids_val = 27'b000000000000000000100000000 ; // (1/128) or 0.00781250
        27'b000010000001000000000000000: neighboring_boids_val = 27'b000000000000000000011111110 ; // (1/129) or 0.00775194
        27'b000010000010000000000000000: neighboring_boids_val = 27'b000000000000000000011111100 ; // (1/130) or 0.00769231
        27'b000010000011000000000000000: neighboring_boids_val = 27'b000000000000000000011111010 ; // (1/131) or 0.00763359
        27'b000010000100000000000000000: neighboring_boids_val = 27'b000000000000000000011111000 ; // (1/132) or 0.00757576
        27'b000010000101000000000000000: neighboring_boids_val = 27'b000000000000000000011110110 ; // (1/133) or 0.00751880
        27'b000010000110000000000000000: neighboring_boids_val = 27'b000000000000000000011110100 ; // (1/134) or 0.00746269
        27'b000010000111000000000000000: neighboring_boids_val = 27'b000000000000000000011110010 ; // (1/135) or 0.00740741
        27'b000010001000000000000000000: neighboring_boids_val = 27'b000000000000000000011110000 ; // (1/136) or 0.00735294
        27'b000010001001000000000000000: neighboring_boids_val = 27'b000000000000000000011101111 ; // (1/137) or 0.00729927
        27'b000010001010000000000000000: neighboring_boids_val = 27'b000000000000000000011101101 ; // (1/138) or 0.00724638
        27'b000010001011000000000000000: neighboring_boids_val = 27'b000000000000000000011101011 ; // (1/139) or 0.00719424
        27'b000010001100000000000000000: neighboring_boids_val = 27'b000000000000000000011101010 ; // (1/140) or 0.00714286
        27'b000010001101000000000000000: neighboring_boids_val = 27'b000000000000000000011101000 ; // (1/141) or 0.00709220
        27'b000010001110000000000000000: neighboring_boids_val = 27'b000000000000000000011100110 ; // (1/142) or 0.00704225
        27'b000010001111000000000000000: neighboring_boids_val = 27'b000000000000000000011100101 ; // (1/143) or 0.00699301
        27'b000010010000000000000000000: neighboring_boids_val = 27'b000000000000000000011100011 ; // (1/144) or 0.00694444
        27'b000010010001000000000000000: neighboring_boids_val = 27'b000000000000000000011100001 ; // (1/145) or 0.00689655
        27'b000010010010000000000000000: neighboring_boids_val = 27'b000000000000000000011100000 ; // (1/146) or 0.00684932
        27'b000010010011000000000000000: neighboring_boids_val = 27'b000000000000000000011011110 ; // (1/147) or 0.00680272
        27'b000010010100000000000000000: neighboring_boids_val = 27'b000000000000000000011011101 ; // (1/148) or 0.00675676
        27'b000010010101000000000000000: neighboring_boids_val = 27'b000000000000000000011011011 ; // (1/149) or 0.00671141
        27'b000010010110000000000000000: neighboring_boids_val = 27'b000000000000000000011011010 ; // (1/150) or 0.00666667
        27'b000010010111000000000000000: neighboring_boids_val = 27'b000000000000000000011011001 ; // (1/151) or 0.00662252
        27'b000010011000000000000000000: neighboring_boids_val = 27'b000000000000000000011010111 ; // (1/152) or 0.00657895
        27'b000010011001000000000000000: neighboring_boids_val = 27'b000000000000000000011010110 ; // (1/153) or 0.00653595
        27'b000010011010000000000000000: neighboring_boids_val = 27'b000000000000000000011010100 ; // (1/154) or 0.00649351
        27'b000010011011000000000000000: neighboring_boids_val = 27'b000000000000000000011010011 ; // (1/155) or 0.00645161
        27'b000010011100000000000000000: neighboring_boids_val = 27'b000000000000000000011010010 ; // (1/156) or 0.00641026
        27'b000010011101000000000000000: neighboring_boids_val = 27'b000000000000000000011010000 ; // (1/157) or 0.00636943
        27'b000010011110000000000000000: neighboring_boids_val = 27'b000000000000000000011001111 ; // (1/158) or 0.00632911
        27'b000010011111000000000000000: neighboring_boids_val = 27'b000000000000000000011001110 ; // (1/159) or 0.00628931
        27'b000010100000000000000000000: neighboring_boids_val = 27'b000000000000000000011001100 ; // (1/160) or 0.00625000
        27'b000010100001000000000000000: neighboring_boids_val = 27'b000000000000000000011001011 ; // (1/161) or 0.00621118
        27'b000010100010000000000000000: neighboring_boids_val = 27'b000000000000000000011001010 ; // (1/162) or 0.00617284
        27'b000010100011000000000000000: neighboring_boids_val = 27'b000000000000000000011001001 ; // (1/163) or 0.00613497
        27'b000010100100000000000000000: neighboring_boids_val = 27'b000000000000000000011000111 ; // (1/164) or 0.00609756
        27'b000010100101000000000000000: neighboring_boids_val = 27'b000000000000000000011000110 ; // (1/165) or 0.00606061
        27'b000010100110000000000000000: neighboring_boids_val = 27'b000000000000000000011000101 ; // (1/166) or 0.00602410
        27'b000010100111000000000000000: neighboring_boids_val = 27'b000000000000000000011000100 ; // (1/167) or 0.00598802
        27'b000010101000000000000000000: neighboring_boids_val = 27'b000000000000000000011000011 ; // (1/168) or 0.00595238
        27'b000010101001000000000000000: neighboring_boids_val = 27'b000000000000000000011000001 ; // (1/169) or 0.00591716
        27'b000010101010000000000000000: neighboring_boids_val = 27'b000000000000000000011000000 ; // (1/170) or 0.00588235
        27'b000010101011000000000000000: neighboring_boids_val = 27'b000000000000000000010111111 ; // (1/171) or 0.00584795
        27'b000010101100000000000000000: neighboring_boids_val = 27'b000000000000000000010111110 ; // (1/172) or 0.00581395
        27'b000010101101000000000000000: neighboring_boids_val = 27'b000000000000000000010111101 ; // (1/173) or 0.00578035
        27'b000010101110000000000000000: neighboring_boids_val = 27'b000000000000000000010111100 ; // (1/174) or 0.00574713
        27'b000010101111000000000000000: neighboring_boids_val = 27'b000000000000000000010111011 ; // (1/175) or 0.00571429
        27'b000010110000000000000000000: neighboring_boids_val = 27'b000000000000000000010111010 ; // (1/176) or 0.00568182
        27'b000010110001000000000000000: neighboring_boids_val = 27'b000000000000000000010111001 ; // (1/177) or 0.00564972
        27'b000010110010000000000000000: neighboring_boids_val = 27'b000000000000000000010111000 ; // (1/178) or 0.00561798
        27'b000010110011000000000000000: neighboring_boids_val = 27'b000000000000000000010110111 ; // (1/179) or 0.00558659
        27'b000010110100000000000000000: neighboring_boids_val = 27'b000000000000000000010110110 ; // (1/180) or 0.00555556
        27'b000010110101000000000000000: neighboring_boids_val = 27'b000000000000000000010110101 ; // (1/181) or 0.00552486
        27'b000010110110000000000000000: neighboring_boids_val = 27'b000000000000000000010110100 ; // (1/182) or 0.00549451
        27'b000010110111000000000000000: neighboring_boids_val = 27'b000000000000000000010110011 ; // (1/183) or 0.00546448
        27'b000010111000000000000000000: neighboring_boids_val = 27'b000000000000000000010110010 ; // (1/184) or 0.00543478
        27'b000010111001000000000000000: neighboring_boids_val = 27'b000000000000000000010110001 ; // (1/185) or 0.00540541
        27'b000010111010000000000000000: neighboring_boids_val = 27'b000000000000000000010110000 ; // (1/186) or 0.00537634
        27'b000010111011000000000000000: neighboring_boids_val = 27'b000000000000000000010101111 ; // (1/187) or 0.00534759
        27'b000010111100000000000000000: neighboring_boids_val = 27'b000000000000000000010101110 ; // (1/188) or 0.00531915
        27'b000010111101000000000000000: neighboring_boids_val = 27'b000000000000000000010101101 ; // (1/189) or 0.00529101
        27'b000010111110000000000000000: neighboring_boids_val = 27'b000000000000000000010101100 ; // (1/190) or 0.00526316
        27'b000010111111000000000000000: neighboring_boids_val = 27'b000000000000000000010101011 ; // (1/191) or 0.00523560
        27'b000011000000000000000000000: neighboring_boids_val = 27'b000000000000000000010101010 ; // (1/192) or 0.00520833
        27'b000011000001000000000000000: neighboring_boids_val = 27'b000000000000000000010101001 ; // (1/193) or 0.00518135
        27'b000011000010000000000000000: neighboring_boids_val = 27'b000000000000000000010101000 ; // (1/194) or 0.00515464
        27'b000011000011000000000000000: neighboring_boids_val = 27'b000000000000000000010101000 ; // (1/195) or 0.00512821
        27'b000011000100000000000000000: neighboring_boids_val = 27'b000000000000000000010100111 ; // (1/196) or 0.00510204
        27'b000011000101000000000000000: neighboring_boids_val = 27'b000000000000000000010100110 ; // (1/197) or 0.00507614
        27'b000011000110000000000000000: neighboring_boids_val = 27'b000000000000000000010100101 ; // (1/198) or 0.00505051
        27'b000011000111000000000000000: neighboring_boids_val = 27'b000000000000000000010100100 ; // (1/199) or 0.00502513
        27'b000011001000000000000000000: neighboring_boids_val = 27'b000000000000000000010100011 ; // (1/200) or 0.00500000
        27'b000011001001000000000000000: neighboring_boids_val = 27'b000000000000000000010100011 ; // (1/201) or 0.00497512
        27'b000011001010000000000000000: neighboring_boids_val = 27'b000000000000000000010100010 ; // (1/202) or 0.00495050
        27'b000011001011000000000000000: neighboring_boids_val = 27'b000000000000000000010100001 ; // (1/203) or 0.00492611
        27'b000011001100000000000000000: neighboring_boids_val = 27'b000000000000000000010100000 ; // (1/204) or 0.00490196
        27'b000011001101000000000000000: neighboring_boids_val = 27'b000000000000000000010011111 ; // (1/205) or 0.00487805
        27'b000011001110000000000000000: neighboring_boids_val = 27'b000000000000000000010011111 ; // (1/206) or 0.00485437
        27'b000011001111000000000000000: neighboring_boids_val = 27'b000000000000000000010011110 ; // (1/207) or 0.00483092
        27'b000011010000000000000000000: neighboring_boids_val = 27'b000000000000000000010011101 ; // (1/208) or 0.00480769
        27'b000011010001000000000000000: neighboring_boids_val = 27'b000000000000000000010011100 ; // (1/209) or 0.00478469
        27'b000011010010000000000000000: neighboring_boids_val = 27'b000000000000000000010011100 ; // (1/210) or 0.00476190
        27'b000011010011000000000000000: neighboring_boids_val = 27'b000000000000000000010011011 ; // (1/211) or 0.00473934
        27'b000011010100000000000000000: neighboring_boids_val = 27'b000000000000000000010011010 ; // (1/212) or 0.00471698
        27'b000011010101000000000000000: neighboring_boids_val = 27'b000000000000000000010011001 ; // (1/213) or 0.00469484
        27'b000011010110000000000000000: neighboring_boids_val = 27'b000000000000000000010011001 ; // (1/214) or 0.00467290
        27'b000011010111000000000000000: neighboring_boids_val = 27'b000000000000000000010011000 ; // (1/215) or 0.00465116
        27'b000011011000000000000000000: neighboring_boids_val = 27'b000000000000000000010010111 ; // (1/216) or 0.00462963
        27'b000011011001000000000000000: neighboring_boids_val = 27'b000000000000000000010010111 ; // (1/217) or 0.00460829
        27'b000011011010000000000000000: neighboring_boids_val = 27'b000000000000000000010010110 ; // (1/218) or 0.00458716
        27'b000011011011000000000000000: neighboring_boids_val = 27'b000000000000000000010010101 ; // (1/219) or 0.00456621
        27'b000011011100000000000000000: neighboring_boids_val = 27'b000000000000000000010010100 ; // (1/220) or 0.00454545
        27'b000011011101000000000000000: neighboring_boids_val = 27'b000000000000000000010010100 ; // (1/221) or 0.00452489
        27'b000011011110000000000000000: neighboring_boids_val = 27'b000000000000000000010010011 ; // (1/222) or 0.00450450
        27'b000011011111000000000000000: neighboring_boids_val = 27'b000000000000000000010010010 ; // (1/223) or 0.00448430
        27'b000011100000000000000000000: neighboring_boids_val = 27'b000000000000000000010010010 ; // (1/224) or 0.00446429
        27'b000011100001000000000000000: neighboring_boids_val = 27'b000000000000000000010010001 ; // (1/225) or 0.00444444
        27'b000011100010000000000000000: neighboring_boids_val = 27'b000000000000000000010010000 ; // (1/226) or 0.00442478
        27'b000011100011000000000000000: neighboring_boids_val = 27'b000000000000000000010010000 ; // (1/227) or 0.00440529
        27'b000011100100000000000000000: neighboring_boids_val = 27'b000000000000000000010001111 ; // (1/228) or 0.00438596
        27'b000011100101000000000000000: neighboring_boids_val = 27'b000000000000000000010001111 ; // (1/229) or 0.00436681
        27'b000011100110000000000000000: neighboring_boids_val = 27'b000000000000000000010001110 ; // (1/230) or 0.00434783
        27'b000011100111000000000000000: neighboring_boids_val = 27'b000000000000000000010001101 ; // (1/231) or 0.00432900
        27'b000011101000000000000000000: neighboring_boids_val = 27'b000000000000000000010001101 ; // (1/232) or 0.00431034
        27'b000011101001000000000000000: neighboring_boids_val = 27'b000000000000000000010001100 ; // (1/233) or 0.00429185
        27'b000011101010000000000000000: neighboring_boids_val = 27'b000000000000000000010001100 ; // (1/234) or 0.00427350
        27'b000011101011000000000000000: neighboring_boids_val = 27'b000000000000000000010001011 ; // (1/235) or 0.00425532
        27'b000011101100000000000000000: neighboring_boids_val = 27'b000000000000000000010001010 ; // (1/236) or 0.00423729
        27'b000011101101000000000000000: neighboring_boids_val = 27'b000000000000000000010001010 ; // (1/237) or 0.00421941
        27'b000011101110000000000000000: neighboring_boids_val = 27'b000000000000000000010001001 ; // (1/238) or 0.00420168
        27'b000011101111000000000000000: neighboring_boids_val = 27'b000000000000000000010001001 ; // (1/239) or 0.00418410
        27'b000011110000000000000000000: neighboring_boids_val = 27'b000000000000000000010001000 ; // (1/240) or 0.00416667
        27'b000011110001000000000000000: neighboring_boids_val = 27'b000000000000000000010000111 ; // (1/241) or 0.00414938
        27'b000011110010000000000000000: neighboring_boids_val = 27'b000000000000000000010000111 ; // (1/242) or 0.00413223
        27'b000011110011000000000000000: neighboring_boids_val = 27'b000000000000000000010000110 ; // (1/243) or 0.00411523
        27'b000011110100000000000000000: neighboring_boids_val = 27'b000000000000000000010000110 ; // (1/244) or 0.00409836
        27'b000011110101000000000000000: neighboring_boids_val = 27'b000000000000000000010000101 ; // (1/245) or 0.00408163
        27'b000011110110000000000000000: neighboring_boids_val = 27'b000000000000000000010000101 ; // (1/246) or 0.00406504
        27'b000011110111000000000000000: neighboring_boids_val = 27'b000000000000000000010000100 ; // (1/247) or 0.00404858
        27'b000011111000000000000000000: neighboring_boids_val = 27'b000000000000000000010000100 ; // (1/248) or 0.00403226
        27'b000011111001000000000000000: neighboring_boids_val = 27'b000000000000000000010000011 ; // (1/249) or 0.00401606
        27'b000011111010000000000000000: neighboring_boids_val = 27'b000000000000000000010000011 ; // (1/250) or 0.00400000
        27'b000011111011000000000000000: neighboring_boids_val = 27'b000000000000000000010000010 ; // (1/251) or 0.00398406
        27'b000011111100000000000000000: neighboring_boids_val = 27'b000000000000000000010000010 ; // (1/252) or 0.00396825
        27'b000011111101000000000000000: neighboring_boids_val = 27'b000000000000000000010000001 ; // (1/253) or 0.00395257
        27'b000011111110000000000000000: neighboring_boids_val = 27'b000000000000000000010000001 ; // (1/254) or 0.00393701
        27'b000011111111000000000000000: neighboring_boids_val = 27'b000000000000000000010000000 ; // (1/255) or 0.00392157
        27'b000100000000000000000000000: neighboring_boids_val = 27'b000000000000000000010000000 ; // (1/256) or 0.00390625
        27'b000100000001000000000000000: neighboring_boids_val = 27'b000000000000000000001111111 ; // (1/257) or 0.00389105
        27'b000100000010000000000000000: neighboring_boids_val = 27'b000000000000000000001111111 ; // (1/258) or 0.00387597
        27'b000100000011000000000000000: neighboring_boids_val = 27'b000000000000000000001111110 ; // (1/259) or 0.00386100
        27'b000100000100000000000000000: neighboring_boids_val = 27'b000000000000000000001111110 ; // (1/260) or 0.00384615
        27'b000100000101000000000000000: neighboring_boids_val = 27'b000000000000000000001111101 ; // (1/261) or 0.00383142
        27'b000100000110000000000000000: neighboring_boids_val = 27'b000000000000000000001111101 ; // (1/262) or 0.00381679
        27'b000100000111000000000000000: neighboring_boids_val = 27'b000000000000000000001111100 ; // (1/263) or 0.00380228
        27'b000100001000000000000000000: neighboring_boids_val = 27'b000000000000000000001111100 ; // (1/264) or 0.00378788
        27'b000100001001000000000000000: neighboring_boids_val = 27'b000000000000000000001111011 ; // (1/265) or 0.00377358
        27'b000100001010000000000000000: neighboring_boids_val = 27'b000000000000000000001111011 ; // (1/266) or 0.00375940
        27'b000100001011000000000000000: neighboring_boids_val = 27'b000000000000000000001111010 ; // (1/267) or 0.00374532
        27'b000100001100000000000000000: neighboring_boids_val = 27'b000000000000000000001111010 ; // (1/268) or 0.00373134
        27'b000100001101000000000000000: neighboring_boids_val = 27'b000000000000000000001111001 ; // (1/269) or 0.00371747
        27'b000100001110000000000000000: neighboring_boids_val = 27'b000000000000000000001111001 ; // (1/270) or 0.00370370
        27'b000100001111000000000000000: neighboring_boids_val = 27'b000000000000000000001111000 ; // (1/271) or 0.00369004
        27'b000100010000000000000000000: neighboring_boids_val = 27'b000000000000000000001111000 ; // (1/272) or 0.00367647
        27'b000100010001000000000000000: neighboring_boids_val = 27'b000000000000000000001111000 ; // (1/273) or 0.00366300
        27'b000100010010000000000000000: neighboring_boids_val = 27'b000000000000000000001110111 ; // (1/274) or 0.00364964
        27'b000100010011000000000000000: neighboring_boids_val = 27'b000000000000000000001110111 ; // (1/275) or 0.00363636
        27'b000100010100000000000000000: neighboring_boids_val = 27'b000000000000000000001110110 ; // (1/276) or 0.00362319
        27'b000100010101000000000000000: neighboring_boids_val = 27'b000000000000000000001110110 ; // (1/277) or 0.00361011
        27'b000100010110000000000000000: neighboring_boids_val = 27'b000000000000000000001110101 ; // (1/278) or 0.00359712
        27'b000100010111000000000000000: neighboring_boids_val = 27'b000000000000000000001110101 ; // (1/279) or 0.00358423
        27'b000100011000000000000000000: neighboring_boids_val = 27'b000000000000000000001110101 ; // (1/280) or 0.00357143
        27'b000100011001000000000000000: neighboring_boids_val = 27'b000000000000000000001110100 ; // (1/281) or 0.00355872
        27'b000100011010000000000000000: neighboring_boids_val = 27'b000000000000000000001110100 ; // (1/282) or 0.00354610
        27'b000100011011000000000000000: neighboring_boids_val = 27'b000000000000000000001110011 ; // (1/283) or 0.00353357
        27'b000100011100000000000000000: neighboring_boids_val = 27'b000000000000000000001110011 ; // (1/284) or 0.00352113
        27'b000100011101000000000000000: neighboring_boids_val = 27'b000000000000000000001110010 ; // (1/285) or 0.00350877
        27'b000100011110000000000000000: neighboring_boids_val = 27'b000000000000000000001110010 ; // (1/286) or 0.00349650
        27'b000100011111000000000000000: neighboring_boids_val = 27'b000000000000000000001110010 ; // (1/287) or 0.00348432
        27'b000100100000000000000000000: neighboring_boids_val = 27'b000000000000000000001110001 ; // (1/288) or 0.00347222
        27'b000100100001000000000000000: neighboring_boids_val = 27'b000000000000000000001110001 ; // (1/289) or 0.00346021
        27'b000100100010000000000000000: neighboring_boids_val = 27'b000000000000000000001110000 ; // (1/290) or 0.00344828
        27'b000100100011000000000000000: neighboring_boids_val = 27'b000000000000000000001110000 ; // (1/291) or 0.00343643
        27'b000100100100000000000000000: neighboring_boids_val = 27'b000000000000000000001110000 ; // (1/292) or 0.00342466
        27'b000100100101000000000000000: neighboring_boids_val = 27'b000000000000000000001101111 ; // (1/293) or 0.00341297
        27'b000100100110000000000000000: neighboring_boids_val = 27'b000000000000000000001101111 ; // (1/294) or 0.00340136
        27'b000100100111000000000000000: neighboring_boids_val = 27'b000000000000000000001101111 ; // (1/295) or 0.00338983
        27'b000100101000000000000000000: neighboring_boids_val = 27'b000000000000000000001101110 ; // (1/296) or 0.00337838
        27'b000100101001000000000000000: neighboring_boids_val = 27'b000000000000000000001101110 ; // (1/297) or 0.00336700
        27'b000100101010000000000000000: neighboring_boids_val = 27'b000000000000000000001101101 ; // (1/298) or 0.00335570
        27'b000100101011000000000000000: neighboring_boids_val = 27'b000000000000000000001101101 ; // (1/299) or 0.00334448
        27'b000100101100000000000000000: neighboring_boids_val = 27'b000000000000000000001101101 ; // (1/300) or 0.00333333
        27'b000100101101000000000000000: neighboring_boids_val = 27'b000000000000000000001101100 ; // (1/301) or 0.00332226
        27'b000100101110000000000000000: neighboring_boids_val = 27'b000000000000000000001101100 ; // (1/302) or 0.00331126
        27'b000100101111000000000000000: neighboring_boids_val = 27'b000000000000000000001101100 ; // (1/303) or 0.00330033
        27'b000100110000000000000000000: neighboring_boids_val = 27'b000000000000000000001101011 ; // (1/304) or 0.00328947
        27'b000100110001000000000000000: neighboring_boids_val = 27'b000000000000000000001101011 ; // (1/305) or 0.00327869
        27'b000100110010000000000000000: neighboring_boids_val = 27'b000000000000000000001101011 ; // (1/306) or 0.00326797
        27'b000100110011000000000000000: neighboring_boids_val = 27'b000000000000000000001101010 ; // (1/307) or 0.00325733
        27'b000100110100000000000000000: neighboring_boids_val = 27'b000000000000000000001101010 ; // (1/308) or 0.00324675
        27'b000100110101000000000000000: neighboring_boids_val = 27'b000000000000000000001101010 ; // (1/309) or 0.00323625
        27'b000100110110000000000000000: neighboring_boids_val = 27'b000000000000000000001101001 ; // (1/310) or 0.00322581
        27'b000100110111000000000000000: neighboring_boids_val = 27'b000000000000000000001101001 ; // (1/311) or 0.00321543
        27'b000100111000000000000000000: neighboring_boids_val = 27'b000000000000000000001101001 ; // (1/312) or 0.00320513
        27'b000100111001000000000000000: neighboring_boids_val = 27'b000000000000000000001101000 ; // (1/313) or 0.00319489
        27'b000100111010000000000000000: neighboring_boids_val = 27'b000000000000000000001101000 ; // (1/314) or 0.00318471
        27'b000100111011000000000000000: neighboring_boids_val = 27'b000000000000000000001101000 ; // (1/315) or 0.00317460
        27'b000100111100000000000000000: neighboring_boids_val = 27'b000000000000000000001100111 ; // (1/316) or 0.00316456
        27'b000100111101000000000000000: neighboring_boids_val = 27'b000000000000000000001100111 ; // (1/317) or 0.00315457
        27'b000100111110000000000000000: neighboring_boids_val = 27'b000000000000000000001100111 ; // (1/318) or 0.00314465
        27'b000100111111000000000000000: neighboring_boids_val = 27'b000000000000000000001100110 ; // (1/319) or 0.00313480
        27'b000101000000000000000000000: neighboring_boids_val = 27'b000000000000000000001100110 ; // (1/320) or 0.00312500
        27'b000101000001000000000000000: neighboring_boids_val = 27'b000000000000000000001100110 ; // (1/321) or 0.00311526
        27'b000101000010000000000000000: neighboring_boids_val = 27'b000000000000000000001100101 ; // (1/322) or 0.00310559
        27'b000101000011000000000000000: neighboring_boids_val = 27'b000000000000000000001100101 ; // (1/323) or 0.00309598
        27'b000101000100000000000000000: neighboring_boids_val = 27'b000000000000000000001100101 ; // (1/324) or 0.00308642
        27'b000101000101000000000000000: neighboring_boids_val = 27'b000000000000000000001100100 ; // (1/325) or 0.00307692
        27'b000101000110000000000000000: neighboring_boids_val = 27'b000000000000000000001100100 ; // (1/326) or 0.00306748
        27'b000101000111000000000000000: neighboring_boids_val = 27'b000000000000000000001100100 ; // (1/327) or 0.00305810
        27'b000101001000000000000000000: neighboring_boids_val = 27'b000000000000000000001100011 ; // (1/328) or 0.00304878
        27'b000101001001000000000000000: neighboring_boids_val = 27'b000000000000000000001100011 ; // (1/329) or 0.00303951
        27'b000101001010000000000000000: neighboring_boids_val = 27'b000000000000000000001100011 ; // (1/330) or 0.00303030
        27'b000101001011000000000000000: neighboring_boids_val = 27'b000000000000000000001100010 ; // (1/331) or 0.00302115
        27'b000101001100000000000000000: neighboring_boids_val = 27'b000000000000000000001100010 ; // (1/332) or 0.00301205
        27'b000101001101000000000000000: neighboring_boids_val = 27'b000000000000000000001100010 ; // (1/333) or 0.00300300
        27'b000101001110000000000000000: neighboring_boids_val = 27'b000000000000000000001100010 ; // (1/334) or 0.00299401
        27'b000101001111000000000000000: neighboring_boids_val = 27'b000000000000000000001100001 ; // (1/335) or 0.00298507
        27'b000101010000000000000000000: neighboring_boids_val = 27'b000000000000000000001100001 ; // (1/336) or 0.00297619
        27'b000101010001000000000000000: neighboring_boids_val = 27'b000000000000000000001100001 ; // (1/337) or 0.00296736
        27'b000101010010000000000000000: neighboring_boids_val = 27'b000000000000000000001100000 ; // (1/338) or 0.00295858
        27'b000101010011000000000000000: neighboring_boids_val = 27'b000000000000000000001100000 ; // (1/339) or 0.00294985
        27'b000101010100000000000000000: neighboring_boids_val = 27'b000000000000000000001100000 ; // (1/340) or 0.00294118
        27'b000101010101000000000000000: neighboring_boids_val = 27'b000000000000000000001100000 ; // (1/341) or 0.00293255
        27'b000101010110000000000000000: neighboring_boids_val = 27'b000000000000000000001011111 ; // (1/342) or 0.00292398
        27'b000101010111000000000000000: neighboring_boids_val = 27'b000000000000000000001011111 ; // (1/343) or 0.00291545
        27'b000101011000000000000000000: neighboring_boids_val = 27'b000000000000000000001011111 ; // (1/344) or 0.00290698
        27'b000101011001000000000000000: neighboring_boids_val = 27'b000000000000000000001011110 ; // (1/345) or 0.00289855
        27'b000101011010000000000000000: neighboring_boids_val = 27'b000000000000000000001011110 ; // (1/346) or 0.00289017
        27'b000101011011000000000000000: neighboring_boids_val = 27'b000000000000000000001011110 ; // (1/347) or 0.00288184
        27'b000101011100000000000000000: neighboring_boids_val = 27'b000000000000000000001011110 ; // (1/348) or 0.00287356
        27'b000101011101000000000000000: neighboring_boids_val = 27'b000000000000000000001011101 ; // (1/349) or 0.00286533
        27'b000101011110000000000000000: neighboring_boids_val = 27'b000000000000000000001011101 ; // (1/350) or 0.00285714
        27'b000101011111000000000000000: neighboring_boids_val = 27'b000000000000000000001011101 ; // (1/351) or 0.00284900
        27'b000101100000000000000000000: neighboring_boids_val = 27'b000000000000000000001011101 ; // (1/352) or 0.00284091
        27'b000101100001000000000000000: neighboring_boids_val = 27'b000000000000000000001011100 ; // (1/353) or 0.00283286
        27'b000101100010000000000000000: neighboring_boids_val = 27'b000000000000000000001011100 ; // (1/354) or 0.00282486
        27'b000101100011000000000000000: neighboring_boids_val = 27'b000000000000000000001011100 ; // (1/355) or 0.00281690
        27'b000101100100000000000000000: neighboring_boids_val = 27'b000000000000000000001011100 ; // (1/356) or 0.00280899
        27'b000101100101000000000000000: neighboring_boids_val = 27'b000000000000000000001011011 ; // (1/357) or 0.00280112
        27'b000101100110000000000000000: neighboring_boids_val = 27'b000000000000000000001011011 ; // (1/358) or 0.00279330
        27'b000101100111000000000000000: neighboring_boids_val = 27'b000000000000000000001011011 ; // (1/359) or 0.00278552
        27'b000101101000000000000000000: neighboring_boids_val = 27'b000000000000000000001011011 ; // (1/360) or 0.00277778
        27'b000101101001000000000000000: neighboring_boids_val = 27'b000000000000000000001011010 ; // (1/361) or 0.00277008
        27'b000101101010000000000000000: neighboring_boids_val = 27'b000000000000000000001011010 ; // (1/362) or 0.00276243
        27'b000101101011000000000000000: neighboring_boids_val = 27'b000000000000000000001011010 ; // (1/363) or 0.00275482
        27'b000101101100000000000000000: neighboring_boids_val = 27'b000000000000000000001011010 ; // (1/364) or 0.00274725
        27'b000101101101000000000000000: neighboring_boids_val = 27'b000000000000000000001011001 ; // (1/365) or 0.00273973
        27'b000101101110000000000000000: neighboring_boids_val = 27'b000000000000000000001011001 ; // (1/366) or 0.00273224
        27'b000101101111000000000000000: neighboring_boids_val = 27'b000000000000000000001011001 ; // (1/367) or 0.00272480
        27'b000101110000000000000000000: neighboring_boids_val = 27'b000000000000000000001011001 ; // (1/368) or 0.00271739
        27'b000101110001000000000000000: neighboring_boids_val = 27'b000000000000000000001011000 ; // (1/369) or 0.00271003
        27'b000101110010000000000000000: neighboring_boids_val = 27'b000000000000000000001011000 ; // (1/370) or 0.00270270
        27'b000101110011000000000000000: neighboring_boids_val = 27'b000000000000000000001011000 ; // (1/371) or 0.00269542
        27'b000101110100000000000000000: neighboring_boids_val = 27'b000000000000000000001011000 ; // (1/372) or 0.00268817
        27'b000101110101000000000000000: neighboring_boids_val = 27'b000000000000000000001010111 ; // (1/373) or 0.00268097
        27'b000101110110000000000000000: neighboring_boids_val = 27'b000000000000000000001010111 ; // (1/374) or 0.00267380
        27'b000101110111000000000000000: neighboring_boids_val = 27'b000000000000000000001010111 ; // (1/375) or 0.00266667
        27'b000101111000000000000000000: neighboring_boids_val = 27'b000000000000000000001010111 ; // (1/376) or 0.00265957
        27'b000101111001000000000000000: neighboring_boids_val = 27'b000000000000000000001010110 ; // (1/377) or 0.00265252
        27'b000101111010000000000000000: neighboring_boids_val = 27'b000000000000000000001010110 ; // (1/378) or 0.00264550
        27'b000101111011000000000000000: neighboring_boids_val = 27'b000000000000000000001010110 ; // (1/379) or 0.00263852
        27'b000101111100000000000000000: neighboring_boids_val = 27'b000000000000000000001010110 ; // (1/380) or 0.00263158
        27'b000101111101000000000000000: neighboring_boids_val = 27'b000000000000000000001010110 ; // (1/381) or 0.00262467
        27'b000101111110000000000000000: neighboring_boids_val = 27'b000000000000000000001010101 ; // (1/382) or 0.00261780
        27'b000101111111000000000000000: neighboring_boids_val = 27'b000000000000000000001010101 ; // (1/383) or 0.00261097
        27'b000110000000000000000000000: neighboring_boids_val = 27'b000000000000000000001010101 ; // (1/384) or 0.00260417
        27'b000110000001000000000000000: neighboring_boids_val = 27'b000000000000000000001010101 ; // (1/385) or 0.00259740
        27'b000110000010000000000000000: neighboring_boids_val = 27'b000000000000000000001010100 ; // (1/386) or 0.00259067
        27'b000110000011000000000000000: neighboring_boids_val = 27'b000000000000000000001010100 ; // (1/387) or 0.00258398
        27'b000110000100000000000000000: neighboring_boids_val = 27'b000000000000000000001010100 ; // (1/388) or 0.00257732
        27'b000110000101000000000000000: neighboring_boids_val = 27'b000000000000000000001010100 ; // (1/389) or 0.00257069
        27'b000110000110000000000000000: neighboring_boids_val = 27'b000000000000000000001010100 ; // (1/390) or 0.00256410
        27'b000110000111000000000000000: neighboring_boids_val = 27'b000000000000000000001010011 ; // (1/391) or 0.00255754
        27'b000110001000000000000000000: neighboring_boids_val = 27'b000000000000000000001010011 ; // (1/392) or 0.00255102
        27'b000110001001000000000000000: neighboring_boids_val = 27'b000000000000000000001010011 ; // (1/393) or 0.00254453
        27'b000110001010000000000000000: neighboring_boids_val = 27'b000000000000000000001010011 ; // (1/394) or 0.00253807
        27'b000110001011000000000000000: neighboring_boids_val = 27'b000000000000000000001010010 ; // (1/395) or 0.00253165
        27'b000110001100000000000000000: neighboring_boids_val = 27'b000000000000000000001010010 ; // (1/396) or 0.00252525
        27'b000110001101000000000000000: neighboring_boids_val = 27'b000000000000000000001010010 ; // (1/397) or 0.00251889
        27'b000110001110000000000000000: neighboring_boids_val = 27'b000000000000000000001010010 ; // (1/398) or 0.00251256
        27'b000110001111000000000000000: neighboring_boids_val = 27'b000000000000000000001010010 ; // (1/399) or 0.00250627
        27'b000110010000000000000000000: neighboring_boids_val = 27'b000000000000000000001010001 ; // (1/400) or 0.00250000
        27'b000110010001000000000000000: neighboring_boids_val = 27'b000000000000000000001010001 ; // (1/401) or 0.00249377
        27'b000110010010000000000000000: neighboring_boids_val = 27'b000000000000000000001010001 ; // (1/402) or 0.00248756
        27'b000110010011000000000000000: neighboring_boids_val = 27'b000000000000000000001010001 ; // (1/403) or 0.00248139
        27'b000110010100000000000000000: neighboring_boids_val = 27'b000000000000000000001010001 ; // (1/404) or 0.00247525
        27'b000110010101000000000000000: neighboring_boids_val = 27'b000000000000000000001010000 ; // (1/405) or 0.00246914
        27'b000110010110000000000000000: neighboring_boids_val = 27'b000000000000000000001010000 ; // (1/406) or 0.00246305
        27'b000110010111000000000000000: neighboring_boids_val = 27'b000000000000000000001010000 ; // (1/407) or 0.00245700
        27'b000110011000000000000000000: neighboring_boids_val = 27'b000000000000000000001010000 ; // (1/408) or 0.00245098
        27'b000110011001000000000000000: neighboring_boids_val = 27'b000000000000000000001010000 ; // (1/409) or 0.00244499
        27'b000110011010000000000000000: neighboring_boids_val = 27'b000000000000000000001001111 ; // (1/410) or 0.00243902
        27'b000110011011000000000000000: neighboring_boids_val = 27'b000000000000000000001001111 ; // (1/411) or 0.00243309
        27'b000110011100000000000000000: neighboring_boids_val = 27'b000000000000000000001001111 ; // (1/412) or 0.00242718
        27'b000110011101000000000000000: neighboring_boids_val = 27'b000000000000000000001001111 ; // (1/413) or 0.00242131
        27'b000110011110000000000000000: neighboring_boids_val = 27'b000000000000000000001001111 ; // (1/414) or 0.00241546
        27'b000110011111000000000000000: neighboring_boids_val = 27'b000000000000000000001001110 ; // (1/415) or 0.00240964
        27'b000110100000000000000000000: neighboring_boids_val = 27'b000000000000000000001001110 ; // (1/416) or 0.00240385
        27'b000110100001000000000000000: neighboring_boids_val = 27'b000000000000000000001001110 ; // (1/417) or 0.00239808
        27'b000110100010000000000000000: neighboring_boids_val = 27'b000000000000000000001001110 ; // (1/418) or 0.00239234
        27'b000110100011000000000000000: neighboring_boids_val = 27'b000000000000000000001001110 ; // (1/419) or 0.00238663
        27'b000110100100000000000000000: neighboring_boids_val = 27'b000000000000000000001001110 ; // (1/420) or 0.00238095
        27'b000110100101000000000000000: neighboring_boids_val = 27'b000000000000000000001001101 ; // (1/421) or 0.00237530
        27'b000110100110000000000000000: neighboring_boids_val = 27'b000000000000000000001001101 ; // (1/422) or 0.00236967
        27'b000110100111000000000000000: neighboring_boids_val = 27'b000000000000000000001001101 ; // (1/423) or 0.00236407
        27'b000110101000000000000000000: neighboring_boids_val = 27'b000000000000000000001001101 ; // (1/424) or 0.00235849
        27'b000110101001000000000000000: neighboring_boids_val = 27'b000000000000000000001001101 ; // (1/425) or 0.00235294
        27'b000110101010000000000000000: neighboring_boids_val = 27'b000000000000000000001001100 ; // (1/426) or 0.00234742
        27'b000110101011000000000000000: neighboring_boids_val = 27'b000000000000000000001001100 ; // (1/427) or 0.00234192
        27'b000110101100000000000000000: neighboring_boids_val = 27'b000000000000000000001001100 ; // (1/428) or 0.00233645
        27'b000110101101000000000000000: neighboring_boids_val = 27'b000000000000000000001001100 ; // (1/429) or 0.00233100
        27'b000110101110000000000000000: neighboring_boids_val = 27'b000000000000000000001001100 ; // (1/430) or 0.00232558
        27'b000110101111000000000000000: neighboring_boids_val = 27'b000000000000000000001001100 ; // (1/431) or 0.00232019
        27'b000110110000000000000000000: neighboring_boids_val = 27'b000000000000000000001001011 ; // (1/432) or 0.00231481
        27'b000110110001000000000000000: neighboring_boids_val = 27'b000000000000000000001001011 ; // (1/433) or 0.00230947
        27'b000110110010000000000000000: neighboring_boids_val = 27'b000000000000000000001001011 ; // (1/434) or 0.00230415
        27'b000110110011000000000000000: neighboring_boids_val = 27'b000000000000000000001001011 ; // (1/435) or 0.00229885
        27'b000110110100000000000000000: neighboring_boids_val = 27'b000000000000000000001001011 ; // (1/436) or 0.00229358
        27'b000110110101000000000000000: neighboring_boids_val = 27'b000000000000000000001001010 ; // (1/437) or 0.00228833
        27'b000110110110000000000000000: neighboring_boids_val = 27'b000000000000000000001001010 ; // (1/438) or 0.00228311
        27'b000110110111000000000000000: neighboring_boids_val = 27'b000000000000000000001001010 ; // (1/439) or 0.00227790
        27'b000110111000000000000000000: neighboring_boids_val = 27'b000000000000000000001001010 ; // (1/440) or 0.00227273
        27'b000110111001000000000000000: neighboring_boids_val = 27'b000000000000000000001001010 ; // (1/441) or 0.00226757
        27'b000110111010000000000000000: neighboring_boids_val = 27'b000000000000000000001001010 ; // (1/442) or 0.00226244
        27'b000110111011000000000000000: neighboring_boids_val = 27'b000000000000000000001001001 ; // (1/443) or 0.00225734
        27'b000110111100000000000000000: neighboring_boids_val = 27'b000000000000000000001001001 ; // (1/444) or 0.00225225
        27'b000110111101000000000000000: neighboring_boids_val = 27'b000000000000000000001001001 ; // (1/445) or 0.00224719
        27'b000110111110000000000000000: neighboring_boids_val = 27'b000000000000000000001001001 ; // (1/446) or 0.00224215
        27'b000110111111000000000000000: neighboring_boids_val = 27'b000000000000000000001001001 ; // (1/447) or 0.00223714
        27'b000111000000000000000000000: neighboring_boids_val = 27'b000000000000000000001001001 ; // (1/448) or 0.00223214
        27'b000111000001000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/449) or 0.00222717
        27'b000111000010000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/450) or 0.00222222
        27'b000111000011000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/451) or 0.00221729
        27'b000111000100000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/452) or 0.00221239
        27'b000111000101000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/453) or 0.00220751
        27'b000111000110000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/454) or 0.00220264
        27'b000111000111000000000000000: neighboring_boids_val = 27'b000000000000000000001001000 ; // (1/455) or 0.00219780
        27'b000111001000000000000000000: neighboring_boids_val = 27'b000000000000000000001000111 ; // (1/456) or 0.00219298
        27'b000111001001000000000000000: neighboring_boids_val = 27'b000000000000000000001000111 ; // (1/457) or 0.00218818
        27'b000111001010000000000000000: neighboring_boids_val = 27'b000000000000000000001000111 ; // (1/458) or 0.00218341
        27'b000111001011000000000000000: neighboring_boids_val = 27'b000000000000000000001000111 ; // (1/459) or 0.00217865
        27'b000111001100000000000000000: neighboring_boids_val = 27'b000000000000000000001000111 ; // (1/460) or 0.00217391
        27'b000111001101000000000000000: neighboring_boids_val = 27'b000000000000000000001000111 ; // (1/461) or 0.00216920
        27'b000111001110000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/462) or 0.00216450
        27'b000111001111000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/463) or 0.00215983
        27'b000111010000000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/464) or 0.00215517
        27'b000111010001000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/465) or 0.00215054
        27'b000111010010000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/466) or 0.00214592
        27'b000111010011000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/467) or 0.00214133
        27'b000111010100000000000000000: neighboring_boids_val = 27'b000000000000000000001000110 ; // (1/468) or 0.00213675
        27'b000111010101000000000000000: neighboring_boids_val = 27'b000000000000000000001000101 ; // (1/469) or 0.00213220
        27'b000111010110000000000000000: neighboring_boids_val = 27'b000000000000000000001000101 ; // (1/470) or 0.00212766
        27'b000111010111000000000000000: neighboring_boids_val = 27'b000000000000000000001000101 ; // (1/471) or 0.00212314
        27'b000111011000000000000000000: neighboring_boids_val = 27'b000000000000000000001000101 ; // (1/472) or 0.00211864
        27'b000111011001000000000000000: neighboring_boids_val = 27'b000000000000000000001000101 ; // (1/473) or 0.00211416
        27'b000111011010000000000000000: neighboring_boids_val = 27'b000000000000000000001000101 ; // (1/474) or 0.00210970
        27'b000111011011000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/475) or 0.00210526
        27'b000111011100000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/476) or 0.00210084
        27'b000111011101000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/477) or 0.00209644
        27'b000111011110000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/478) or 0.00209205
        27'b000111011111000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/479) or 0.00208768
        27'b000111100000000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/480) or 0.00208333
        27'b000111100001000000000000000: neighboring_boids_val = 27'b000000000000000000001000100 ; // (1/481) or 0.00207900
        27'b000111100010000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/482) or 0.00207469
        27'b000111100011000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/483) or 0.00207039
        27'b000111100100000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/484) or 0.00206612
        27'b000111100101000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/485) or 0.00206186
        27'b000111100110000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/486) or 0.00205761
        27'b000111100111000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/487) or 0.00205339
        27'b000111101000000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/488) or 0.00204918
        27'b000111101001000000000000000: neighboring_boids_val = 27'b000000000000000000001000011 ; // (1/489) or 0.00204499
        27'b000111101010000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/490) or 0.00204082
        27'b000111101011000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/491) or 0.00203666
        27'b000111101100000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/492) or 0.00203252
        27'b000111101101000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/493) or 0.00202840
        27'b000111101110000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/494) or 0.00202429
        27'b000111101111000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/495) or 0.00202020
        27'b000111110000000000000000000: neighboring_boids_val = 27'b000000000000000000001000010 ; // (1/496) or 0.00201613
        27'b000111110001000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/497) or 0.00201207
        27'b000111110010000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/498) or 0.00200803
        27'b000111110011000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/499) or 0.00200401
        27'b000111110100000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/500) or 0.00200000
        27'b000111110101000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/501) or 0.00199601
        27'b000111110110000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/502) or 0.00199203
        27'b000111110111000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/503) or 0.00198807
        27'b000111111000000000000000000: neighboring_boids_val = 27'b000000000000000000001000001 ; // (1/504) or 0.00198413
        27'b000111111001000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/505) or 0.00198020
        27'b000111111010000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/506) or 0.00197628
        27'b000111111011000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/507) or 0.00197239
        27'b000111111100000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/508) or 0.00196850
        27'b000111111101000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/509) or 0.00196464
        27'b000111111110000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/510) or 0.00196078
        27'b000111111111000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/511) or 0.00195695
        27'b001000000000000000000000000: neighboring_boids_val = 27'b000000000000000000001000000 ; // (1/512) or 0.00195312
        27'b001000000001000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/513) or 0.00194932
        27'b001000000010000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/514) or 0.00194553
        27'b001000000011000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/515) or 0.00194175
        27'b001000000100000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/516) or 0.00193798
        27'b001000000101000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/517) or 0.00193424
        27'b001000000110000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/518) or 0.00193050
        27'b001000000111000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/519) or 0.00192678
        27'b001000001000000000000000000: neighboring_boids_val = 27'b000000000000000000000111111 ; // (1/520) or 0.00192308
        27'b001000001001000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/521) or 0.00191939
        27'b001000001010000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/522) or 0.00191571
        27'b001000001011000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/523) or 0.00191205
        27'b001000001100000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/524) or 0.00190840
        27'b001000001101000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/525) or 0.00190476
        27'b001000001110000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/526) or 0.00190114
        27'b001000001111000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/527) or 0.00189753
        27'b001000010000000000000000000: neighboring_boids_val = 27'b000000000000000000000111110 ; // (1/528) or 0.00189394
        27'b001000010001000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/529) or 0.00189036
        27'b001000010010000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/530) or 0.00188679
        27'b001000010011000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/531) or 0.00188324
        27'b001000010100000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/532) or 0.00187970
        27'b001000010101000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/533) or 0.00187617
        27'b001000010110000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/534) or 0.00187266
        27'b001000010111000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/535) or 0.00186916
        27'b001000011000000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/536) or 0.00186567
        27'b001000011001000000000000000: neighboring_boids_val = 27'b000000000000000000000111101 ; // (1/537) or 0.00186220
        27'b001000011010000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/538) or 0.00185874
        27'b001000011011000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/539) or 0.00185529
        27'b001000011100000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/540) or 0.00185185
        27'b001000011101000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/541) or 0.00184843
        27'b001000011110000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/542) or 0.00184502
        27'b001000011111000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/543) or 0.00184162
        27'b001000100000000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/544) or 0.00183824
        27'b001000100001000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/545) or 0.00183486
        27'b001000100010000000000000000: neighboring_boids_val = 27'b000000000000000000000111100 ; // (1/546) or 0.00183150
        27'b001000100011000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/547) or 0.00182815
        27'b001000100100000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/548) or 0.00182482
        27'b001000100101000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/549) or 0.00182149
        27'b001000100110000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/550) or 0.00181818
        27'b001000100111000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/551) or 0.00181488
        27'b001000101000000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/552) or 0.00181159
        27'b001000101001000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/553) or 0.00180832
        27'b001000101010000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/554) or 0.00180505
        27'b001000101011000000000000000: neighboring_boids_val = 27'b000000000000000000000111011 ; // (1/555) or 0.00180180
        27'b001000101100000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/556) or 0.00179856
        27'b001000101101000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/557) or 0.00179533
        27'b001000101110000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/558) or 0.00179211
        27'b001000101111000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/559) or 0.00178891
        27'b001000110000000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/560) or 0.00178571
        27'b001000110001000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/561) or 0.00178253
        27'b001000110010000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/562) or 0.00177936
        27'b001000110011000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/563) or 0.00177620
        27'b001000110100000000000000000: neighboring_boids_val = 27'b000000000000000000000111010 ; // (1/564) or 0.00177305
        27'b001000110101000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/565) or 0.00176991
        27'b001000110110000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/566) or 0.00176678
        27'b001000110111000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/567) or 0.00176367
        27'b001000111000000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/568) or 0.00176056
        27'b001000111001000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/569) or 0.00175747
        27'b001000111010000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/570) or 0.00175439
        27'b001000111011000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/571) or 0.00175131
        27'b001000111100000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/572) or 0.00174825
        27'b001000111101000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/573) or 0.00174520
        27'b001000111110000000000000000: neighboring_boids_val = 27'b000000000000000000000111001 ; // (1/574) or 0.00174216
        27'b001000111111000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/575) or 0.00173913
        27'b001001000000000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/576) or 0.00173611
        27'b001001000001000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/577) or 0.00173310
        27'b001001000010000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/578) or 0.00173010
        27'b001001000011000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/579) or 0.00172712
        27'b001001000100000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/580) or 0.00172414
        27'b001001000101000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/581) or 0.00172117
        27'b001001000110000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/582) or 0.00171821
        27'b001001000111000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/583) or 0.00171527
        27'b001001001000000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/584) or 0.00171233
        27'b001001001001000000000000000: neighboring_boids_val = 27'b000000000000000000000111000 ; // (1/585) or 0.00170940
        27'b001001001010000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/586) or 0.00170648
        27'b001001001011000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/587) or 0.00170358
        27'b001001001100000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/588) or 0.00170068
        27'b001001001101000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/589) or 0.00169779
        27'b001001001110000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/590) or 0.00169492
        27'b001001001111000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/591) or 0.00169205
        27'b001001010000000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/592) or 0.00168919
        27'b001001010001000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/593) or 0.00168634
        27'b001001010010000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/594) or 0.00168350
        27'b001001010011000000000000000: neighboring_boids_val = 27'b000000000000000000000110111 ; // (1/595) or 0.00168067
        27'b001001010100000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/596) or 0.00167785
        27'b001001010101000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/597) or 0.00167504
        27'b001001010110000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/598) or 0.00167224
        27'b001001010111000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/599) or 0.00166945
        27'b001001011000000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/600) or 0.00166667
        27'b001001011001000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/601) or 0.00166389
        27'b001001011010000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/602) or 0.00166113
        27'b001001011011000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/603) or 0.00165837
        27'b001001011100000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/604) or 0.00165563
        27'b001001011101000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/605) or 0.00165289
        27'b001001011110000000000000000: neighboring_boids_val = 27'b000000000000000000000110110 ; // (1/606) or 0.00165017
        27'b001001011111000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/607) or 0.00164745
        27'b001001100000000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/608) or 0.00164474
        27'b001001100001000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/609) or 0.00164204
        27'b001001100010000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/610) or 0.00163934
        27'b001001100011000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/611) or 0.00163666
        27'b001001100100000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/612) or 0.00163399
        27'b001001100101000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/613) or 0.00163132
        27'b001001100110000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/614) or 0.00162866
        27'b001001100111000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/615) or 0.00162602
        27'b001001101000000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/616) or 0.00162338
        27'b001001101001000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/617) or 0.00162075
        27'b001001101010000000000000000: neighboring_boids_val = 27'b000000000000000000000110101 ; // (1/618) or 0.00161812
        27'b001001101011000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/619) or 0.00161551
        27'b001001101100000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/620) or 0.00161290
        27'b001001101101000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/621) or 0.00161031
        27'b001001101110000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/622) or 0.00160772
        27'b001001101111000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/623) or 0.00160514
        27'b001001110000000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/624) or 0.00160256
        27'b001001110001000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/625) or 0.00160000
        27'b001001110010000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/626) or 0.00159744
        27'b001001110011000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/627) or 0.00159490
        27'b001001110100000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/628) or 0.00159236
        27'b001001110101000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/629) or 0.00158983
        27'b001001110110000000000000000: neighboring_boids_val = 27'b000000000000000000000110100 ; // (1/630) or 0.00158730
        27'b001001110111000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/631) or 0.00158479
        27'b001001111000000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/632) or 0.00158228
        27'b001001111001000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/633) or 0.00157978
        27'b001001111010000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/634) or 0.00157729
        27'b001001111011000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/635) or 0.00157480
        27'b001001111100000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/636) or 0.00157233
        27'b001001111101000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/637) or 0.00156986
        27'b001001111110000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/638) or 0.00156740
        27'b001001111111000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/639) or 0.00156495
        27'b001010000000000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/640) or 0.00156250
        27'b001010000001000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/641) or 0.00156006
        27'b001010000010000000000000000: neighboring_boids_val = 27'b000000000000000000000110011 ; // (1/642) or 0.00155763
        27'b001010000011000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/643) or 0.00155521
        27'b001010000100000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/644) or 0.00155280
        27'b001010000101000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/645) or 0.00155039
        27'b001010000110000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/646) or 0.00154799
        27'b001010000111000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/647) or 0.00154560
        27'b001010001000000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/648) or 0.00154321
        27'b001010001001000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/649) or 0.00154083
        27'b001010001010000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/650) or 0.00153846
        27'b001010001011000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/651) or 0.00153610
        27'b001010001100000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/652) or 0.00153374
        27'b001010001101000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/653) or 0.00153139
        27'b001010001110000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/654) or 0.00152905
        27'b001010001111000000000000000: neighboring_boids_val = 27'b000000000000000000000110010 ; // (1/655) or 0.00152672
        27'b001010010000000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/656) or 0.00152439
        27'b001010010001000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/657) or 0.00152207
        27'b001010010010000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/658) or 0.00151976
        27'b001010010011000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/659) or 0.00151745
        27'b001010010100000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/660) or 0.00151515
        27'b001010010101000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/661) or 0.00151286
        27'b001010010110000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/662) or 0.00151057
        27'b001010010111000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/663) or 0.00150830
        27'b001010011000000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/664) or 0.00150602
        27'b001010011001000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/665) or 0.00150376
        27'b001010011010000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/666) or 0.00150150
        27'b001010011011000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/667) or 0.00149925
        27'b001010011100000000000000000: neighboring_boids_val = 27'b000000000000000000000110001 ; // (1/668) or 0.00149701
        27'b001010011101000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/669) or 0.00149477
        27'b001010011110000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/670) or 0.00149254
        27'b001010011111000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/671) or 0.00149031
        27'b001010100000000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/672) or 0.00148810
        27'b001010100001000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/673) or 0.00148588
        27'b001010100010000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/674) or 0.00148368
        27'b001010100011000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/675) or 0.00148148
        27'b001010100100000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/676) or 0.00147929
        27'b001010100101000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/677) or 0.00147710
        27'b001010100110000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/678) or 0.00147493
        27'b001010100111000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/679) or 0.00147275
        27'b001010101000000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/680) or 0.00147059
        27'b001010101001000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/681) or 0.00146843
        27'b001010101010000000000000000: neighboring_boids_val = 27'b000000000000000000000110000 ; // (1/682) or 0.00146628
        27'b001010101011000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/683) or 0.00146413
        27'b001010101100000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/684) or 0.00146199
        27'b001010101101000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/685) or 0.00145985
        27'b001010101110000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/686) or 0.00145773
        27'b001010101111000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/687) or 0.00145560
        27'b001010110000000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/688) or 0.00145349
        27'b001010110001000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/689) or 0.00145138
        27'b001010110010000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/690) or 0.00144928
        27'b001010110011000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/691) or 0.00144718
        27'b001010110100000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/692) or 0.00144509
        27'b001010110101000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/693) or 0.00144300
        27'b001010110110000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/694) or 0.00144092
        27'b001010110111000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/695) or 0.00143885
        27'b001010111000000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/696) or 0.00143678
        27'b001010111001000000000000000: neighboring_boids_val = 27'b000000000000000000000101111 ; // (1/697) or 0.00143472
        27'b001010111010000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/698) or 0.00143266
        27'b001010111011000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/699) or 0.00143062
        27'b001010111100000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/700) or 0.00142857
        27'b001010111101000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/701) or 0.00142653
        27'b001010111110000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/702) or 0.00142450
        27'b001010111111000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/703) or 0.00142248
        27'b001011000000000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/704) or 0.00142045
        27'b001011000001000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/705) or 0.00141844
        27'b001011000010000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/706) or 0.00141643
        27'b001011000011000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/707) or 0.00141443
        27'b001011000100000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/708) or 0.00141243
        27'b001011000101000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/709) or 0.00141044
        27'b001011000110000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/710) or 0.00140845
        27'b001011000111000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/711) or 0.00140647
        27'b001011001000000000000000000: neighboring_boids_val = 27'b000000000000000000000101110 ; // (1/712) or 0.00140449
        27'b001011001001000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/713) or 0.00140252
        27'b001011001010000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/714) or 0.00140056
        27'b001011001011000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/715) or 0.00139860
        27'b001011001100000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/716) or 0.00139665
        27'b001011001101000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/717) or 0.00139470
        27'b001011001110000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/718) or 0.00139276
        27'b001011001111000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/719) or 0.00139082
        27'b001011010000000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/720) or 0.00138889
        27'b001011010001000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/721) or 0.00138696
        27'b001011010010000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/722) or 0.00138504
        27'b001011010011000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/723) or 0.00138313
        27'b001011010100000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/724) or 0.00138122
        27'b001011010101000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/725) or 0.00137931
        27'b001011010110000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/726) or 0.00137741
        27'b001011010111000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/727) or 0.00137552
        27'b001011011000000000000000000: neighboring_boids_val = 27'b000000000000000000000101101 ; // (1/728) or 0.00137363
        27'b001011011001000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/729) or 0.00137174
        27'b001011011010000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/730) or 0.00136986
        27'b001011011011000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/731) or 0.00136799
        27'b001011011100000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/732) or 0.00136612
        27'b001011011101000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/733) or 0.00136426
        27'b001011011110000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/734) or 0.00136240
        27'b001011011111000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/735) or 0.00136054
        27'b001011100000000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/736) or 0.00135870
        27'b001011100001000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/737) or 0.00135685
        27'b001011100010000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/738) or 0.00135501
        27'b001011100011000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/739) or 0.00135318
        27'b001011100100000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/740) or 0.00135135
        27'b001011100101000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/741) or 0.00134953
        27'b001011100110000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/742) or 0.00134771
        27'b001011100111000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/743) or 0.00134590
        27'b001011101000000000000000000: neighboring_boids_val = 27'b000000000000000000000101100 ; // (1/744) or 0.00134409
        27'b001011101001000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/745) or 0.00134228
        27'b001011101010000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/746) or 0.00134048
        27'b001011101011000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/747) or 0.00133869
        27'b001011101100000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/748) or 0.00133690
        27'b001011101101000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/749) or 0.00133511
        27'b001011101110000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/750) or 0.00133333
        27'b001011101111000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/751) or 0.00133156
        27'b001011110000000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/752) or 0.00132979
        27'b001011110001000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/753) or 0.00132802
        27'b001011110010000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/754) or 0.00132626
        27'b001011110011000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/755) or 0.00132450
        27'b001011110100000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/756) or 0.00132275
        27'b001011110101000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/757) or 0.00132100
        27'b001011110110000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/758) or 0.00131926
        27'b001011110111000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/759) or 0.00131752
        27'b001011111000000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/760) or 0.00131579
        27'b001011111001000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/761) or 0.00131406
        27'b001011111010000000000000000: neighboring_boids_val = 27'b000000000000000000000101011 ; // (1/762) or 0.00131234
        27'b001011111011000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/763) or 0.00131062
        27'b001011111100000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/764) or 0.00130890
        27'b001011111101000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/765) or 0.00130719
        27'b001011111110000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/766) or 0.00130548
        27'b001011111111000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/767) or 0.00130378
        27'b001100000000000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/768) or 0.00130208
        27'b001100000001000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/769) or 0.00130039
        27'b001100000010000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/770) or 0.00129870
        27'b001100000011000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/771) or 0.00129702
        27'b001100000100000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/772) or 0.00129534
        27'b001100000101000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/773) or 0.00129366
        27'b001100000110000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/774) or 0.00129199
        27'b001100000111000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/775) or 0.00129032
        27'b001100001000000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/776) or 0.00128866
        27'b001100001001000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/777) or 0.00128700
        27'b001100001010000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/778) or 0.00128535
        27'b001100001011000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/779) or 0.00128370
        27'b001100001100000000000000000: neighboring_boids_val = 27'b000000000000000000000101010 ; // (1/780) or 0.00128205
        27'b001100001101000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/781) or 0.00128041
        27'b001100001110000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/782) or 0.00127877
        27'b001100001111000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/783) or 0.00127714
        27'b001100010000000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/784) or 0.00127551
        27'b001100010001000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/785) or 0.00127389
        27'b001100010010000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/786) or 0.00127226
        27'b001100010011000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/787) or 0.00127065
        27'b001100010100000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/788) or 0.00126904
        27'b001100010101000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/789) or 0.00126743
        27'b001100010110000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/790) or 0.00126582
        27'b001100010111000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/791) or 0.00126422
        27'b001100011000000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/792) or 0.00126263
        27'b001100011001000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/793) or 0.00126103
        27'b001100011010000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/794) or 0.00125945
        27'b001100011011000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/795) or 0.00125786
        27'b001100011100000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/796) or 0.00125628
        27'b001100011101000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/797) or 0.00125471
        27'b001100011110000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/798) or 0.00125313
        27'b001100011111000000000000000: neighboring_boids_val = 27'b000000000000000000000101001 ; // (1/799) or 0.00125156
        27'b001100100000000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/800) or 0.00125000
        27'b001100100001000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/801) or 0.00124844
        27'b001100100010000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/802) or 0.00124688
        27'b001100100011000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/803) or 0.00124533
        27'b001100100100000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/804) or 0.00124378
        27'b001100100101000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/805) or 0.00124224
        27'b001100100110000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/806) or 0.00124069
        27'b001100100111000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/807) or 0.00123916
        27'b001100101000000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/808) or 0.00123762
        27'b001100101001000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/809) or 0.00123609
        27'b001100101010000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/810) or 0.00123457
        27'b001100101011000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/811) or 0.00123305
        27'b001100101100000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/812) or 0.00123153
        27'b001100101101000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/813) or 0.00123001
        27'b001100101110000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/814) or 0.00122850
        27'b001100101111000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/815) or 0.00122699
        27'b001100110000000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/816) or 0.00122549
        27'b001100110001000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/817) or 0.00122399
        27'b001100110010000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/818) or 0.00122249
        27'b001100110011000000000000000: neighboring_boids_val = 27'b000000000000000000000101000 ; // (1/819) or 0.00122100
        27'b001100110100000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/820) or 0.00121951
        27'b001100110101000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/821) or 0.00121803
        27'b001100110110000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/822) or 0.00121655
        27'b001100110111000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/823) or 0.00121507
        27'b001100111000000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/824) or 0.00121359
        27'b001100111001000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/825) or 0.00121212
        27'b001100111010000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/826) or 0.00121065
        27'b001100111011000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/827) or 0.00120919
        27'b001100111100000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/828) or 0.00120773
        27'b001100111101000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/829) or 0.00120627
        27'b001100111110000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/830) or 0.00120482
        27'b001100111111000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/831) or 0.00120337
        27'b001101000000000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/832) or 0.00120192
        27'b001101000001000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/833) or 0.00120048
        27'b001101000010000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/834) or 0.00119904
        27'b001101000011000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/835) or 0.00119760
        27'b001101000100000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/836) or 0.00119617
        27'b001101000101000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/837) or 0.00119474
        27'b001101000110000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/838) or 0.00119332
        27'b001101000111000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/839) or 0.00119190
        27'b001101001000000000000000000: neighboring_boids_val = 27'b000000000000000000000100111 ; // (1/840) or 0.00119048
        27'b001101001001000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/841) or 0.00118906
        27'b001101001010000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/842) or 0.00118765
        27'b001101001011000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/843) or 0.00118624
        27'b001101001100000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/844) or 0.00118483
        27'b001101001101000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/845) or 0.00118343
        27'b001101001110000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/846) or 0.00118203
        27'b001101001111000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/847) or 0.00118064
        27'b001101010000000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/848) or 0.00117925
        27'b001101010001000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/849) or 0.00117786
        27'b001101010010000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/850) or 0.00117647
        27'b001101010011000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/851) or 0.00117509
        27'b001101010100000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/852) or 0.00117371
        27'b001101010101000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/853) or 0.00117233
        27'b001101010110000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/854) or 0.00117096
        27'b001101010111000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/855) or 0.00116959
        27'b001101011000000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/856) or 0.00116822
        27'b001101011001000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/857) or 0.00116686
        27'b001101011010000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/858) or 0.00116550
        27'b001101011011000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/859) or 0.00116414
        27'b001101011100000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/860) or 0.00116279
        27'b001101011101000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/861) or 0.00116144
        27'b001101011110000000000000000: neighboring_boids_val = 27'b000000000000000000000100110 ; // (1/862) or 0.00116009
        27'b001101011111000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/863) or 0.00115875
        27'b001101100000000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/864) or 0.00115741
        27'b001101100001000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/865) or 0.00115607
        27'b001101100010000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/866) or 0.00115473
        27'b001101100011000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/867) or 0.00115340
        27'b001101100100000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/868) or 0.00115207
        27'b001101100101000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/869) or 0.00115075
        27'b001101100110000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/870) or 0.00114943
        27'b001101100111000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/871) or 0.00114811
        27'b001101101000000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/872) or 0.00114679
        27'b001101101001000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/873) or 0.00114548
        27'b001101101010000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/874) or 0.00114416
        27'b001101101011000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/875) or 0.00114286
        27'b001101101100000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/876) or 0.00114155
        27'b001101101101000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/877) or 0.00114025
        27'b001101101110000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/878) or 0.00113895
        27'b001101101111000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/879) or 0.00113766
        27'b001101110000000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/880) or 0.00113636
        27'b001101110001000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/881) or 0.00113507
        27'b001101110010000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/882) or 0.00113379
        27'b001101110011000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/883) or 0.00113250
        27'b001101110100000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/884) or 0.00113122
        27'b001101110101000000000000000: neighboring_boids_val = 27'b000000000000000000000100101 ; // (1/885) or 0.00112994
        27'b001101110110000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/886) or 0.00112867
        27'b001101110111000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/887) or 0.00112740
        27'b001101111000000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/888) or 0.00112613
        27'b001101111001000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/889) or 0.00112486
        27'b001101111010000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/890) or 0.00112360
        27'b001101111011000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/891) or 0.00112233
        27'b001101111100000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/892) or 0.00112108
        27'b001101111101000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/893) or 0.00111982
        27'b001101111110000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/894) or 0.00111857
        27'b001101111111000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/895) or 0.00111732
        27'b001110000000000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/896) or 0.00111607
        27'b001110000001000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/897) or 0.00111483
        27'b001110000010000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/898) or 0.00111359
        27'b001110000011000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/899) or 0.00111235
        27'b001110000100000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/900) or 0.00111111
        27'b001110000101000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/901) or 0.00110988
        27'b001110000110000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/902) or 0.00110865
        27'b001110000111000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/903) or 0.00110742
        27'b001110001000000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/904) or 0.00110619
        27'b001110001001000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/905) or 0.00110497
        27'b001110001010000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/906) or 0.00110375
        27'b001110001011000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/907) or 0.00110254
        27'b001110001100000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/908) or 0.00110132
        27'b001110001101000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/909) or 0.00110011
        27'b001110001110000000000000000: neighboring_boids_val = 27'b000000000000000000000100100 ; // (1/910) or 0.00109890
        27'b001110001111000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/911) or 0.00109769
        27'b001110010000000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/912) or 0.00109649
        27'b001110010001000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/913) or 0.00109529
        27'b001110010010000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/914) or 0.00109409
        27'b001110010011000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/915) or 0.00109290
        27'b001110010100000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/916) or 0.00109170
        27'b001110010101000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/917) or 0.00109051
        27'b001110010110000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/918) or 0.00108932
        27'b001110010111000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/919) or 0.00108814
        27'b001110011000000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/920) or 0.00108696
        27'b001110011001000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/921) or 0.00108578
        27'b001110011010000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/922) or 0.00108460
        27'b001110011011000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/923) or 0.00108342
        27'b001110011100000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/924) or 0.00108225
        27'b001110011101000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/925) or 0.00108108
        27'b001110011110000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/926) or 0.00107991
        27'b001110011111000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/927) or 0.00107875
        27'b001110100000000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/928) or 0.00107759
        27'b001110100001000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/929) or 0.00107643
        27'b001110100010000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/930) or 0.00107527
        27'b001110100011000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/931) or 0.00107411
        27'b001110100100000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/932) or 0.00107296
        27'b001110100101000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/933) or 0.00107181
        27'b001110100110000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/934) or 0.00107066
        27'b001110100111000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/935) or 0.00106952
        27'b001110101000000000000000000: neighboring_boids_val = 27'b000000000000000000000100011 ; // (1/936) or 0.00106838
        27'b001110101001000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/937) or 0.00106724
        27'b001110101010000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/938) or 0.00106610
        27'b001110101011000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/939) or 0.00106496
        27'b001110101100000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/940) or 0.00106383
        27'b001110101101000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/941) or 0.00106270
        27'b001110101110000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/942) or 0.00106157
        27'b001110101111000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/943) or 0.00106045
        27'b001110110000000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/944) or 0.00105932
        27'b001110110001000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/945) or 0.00105820
        27'b001110110010000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/946) or 0.00105708
        27'b001110110011000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/947) or 0.00105597
        27'b001110110100000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/948) or 0.00105485
        27'b001110110101000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/949) or 0.00105374
        27'b001110110110000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/950) or 0.00105263
        27'b001110110111000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/951) or 0.00105152
        27'b001110111000000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/952) or 0.00105042
        27'b001110111001000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/953) or 0.00104932
        27'b001110111010000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/954) or 0.00104822
        27'b001110111011000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/955) or 0.00104712
        27'b001110111100000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/956) or 0.00104603
        27'b001110111101000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/957) or 0.00104493
        27'b001110111110000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/958) or 0.00104384
        27'b001110111111000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/959) or 0.00104275
        27'b001111000000000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/960) or 0.00104167
        27'b001111000001000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/961) or 0.00104058
        27'b001111000010000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/962) or 0.00103950
        27'b001111000011000000000000000: neighboring_boids_val = 27'b000000000000000000000100010 ; // (1/963) or 0.00103842
        27'b001111000100000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/964) or 0.00103734
        27'b001111000101000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/965) or 0.00103627
        27'b001111000110000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/966) or 0.00103520
        27'b001111000111000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/967) or 0.00103413
        27'b001111001000000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/968) or 0.00103306
        27'b001111001001000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/969) or 0.00103199
        27'b001111001010000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/970) or 0.00103093
        27'b001111001011000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/971) or 0.00102987
        27'b001111001100000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/972) or 0.00102881
        27'b001111001101000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/973) or 0.00102775
        27'b001111001110000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/974) or 0.00102669
        27'b001111001111000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/975) or 0.00102564
        27'b001111010000000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/976) or 0.00102459
        27'b001111010001000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/977) or 0.00102354
        27'b001111010010000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/978) or 0.00102249
        27'b001111010011000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/979) or 0.00102145
        27'b001111010100000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/980) or 0.00102041
        27'b001111010101000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/981) or 0.00101937
        27'b001111010110000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/982) or 0.00101833
        27'b001111010111000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/983) or 0.00101729
        27'b001111011000000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/984) or 0.00101626
        27'b001111011001000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/985) or 0.00101523
        27'b001111011010000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/986) or 0.00101420
        27'b001111011011000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/987) or 0.00101317
        27'b001111011100000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/988) or 0.00101215
        27'b001111011101000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/989) or 0.00101112
        27'b001111011110000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/990) or 0.00101010
        27'b001111011111000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/991) or 0.00100908
        27'b001111100000000000000000000: neighboring_boids_val = 27'b000000000000000000000100001 ; // (1/992) or 0.00100806
        27'b001111100001000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/993) or 0.00100705
        27'b001111100010000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/994) or 0.00100604
        27'b001111100011000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/995) or 0.00100503
        27'b001111100100000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/996) or 0.00100402
        27'b001111100101000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/997) or 0.00100301
        27'b001111100110000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/998) or 0.00100200
        27'b001111100111000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/999) or 0.00100100
        27'b001111101000000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1000) or 0.00100000
        27'b001111101001000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1001) or 0.00099900
        27'b001111101010000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1002) or 0.00099800
        27'b001111101011000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1003) or 0.00099701
        27'b001111101100000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1004) or 0.00099602
        27'b001111101101000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1005) or 0.00099502
        27'b001111101110000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1006) or 0.00099404
        27'b001111101111000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1007) or 0.00099305
        27'b001111110000000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1008) or 0.00099206
        27'b001111110001000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1009) or 0.00099108
        27'b001111110010000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1010) or 0.00099010
        27'b001111110011000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1011) or 0.00098912
        27'b001111110100000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1012) or 0.00098814
        27'b001111110101000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1013) or 0.00098717
        27'b001111110110000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1014) or 0.00098619
        27'b001111110111000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1015) or 0.00098522
        27'b001111111000000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1016) or 0.00098425
        27'b001111111001000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1017) or 0.00098328
        27'b001111111010000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1018) or 0.00098232
        27'b001111111011000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1019) or 0.00098135
        27'b001111111100000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1020) or 0.00098039
        27'b001111111101000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1021) or 0.00097943
        27'b001111111110000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1022) or 0.00097847
        27'b001111111111000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1023) or 0.00097752
        27'b010000000000000000000000000: neighboring_boids_val = 27'b000000000000000000000100000 ; // (1/1024) or 0.00097656
        27'b010000000001000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1025) or 0.00097561
        27'b010000000010000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1026) or 0.00097466
        27'b010000000011000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1027) or 0.00097371
        27'b010000000100000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1028) or 0.00097276
        27'b010000000101000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1029) or 0.00097182
        27'b010000000110000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1030) or 0.00097087
        27'b010000000111000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1031) or 0.00096993
        27'b010000001000000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1032) or 0.00096899
        27'b010000001001000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1033) or 0.00096805
        27'b010000001010000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1034) or 0.00096712
        27'b010000001011000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1035) or 0.00096618
        27'b010000001100000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1036) or 0.00096525
        27'b010000001101000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1037) or 0.00096432
        27'b010000001110000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1038) or 0.00096339
        27'b010000001111000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1039) or 0.00096246
        27'b010000010000000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1040) or 0.00096154
        27'b010000010001000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1041) or 0.00096061
        27'b010000010010000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1042) or 0.00095969
        27'b010000010011000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1043) or 0.00095877
        27'b010000010100000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1044) or 0.00095785
        27'b010000010101000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1045) or 0.00095694
        27'b010000010110000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1046) or 0.00095602
        27'b010000010111000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1047) or 0.00095511
        27'b010000011000000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1048) or 0.00095420
        27'b010000011001000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1049) or 0.00095329
        27'b010000011010000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1050) or 0.00095238
        27'b010000011011000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1051) or 0.00095147
        27'b010000011100000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1052) or 0.00095057
        27'b010000011101000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1053) or 0.00094967
        27'b010000011110000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1054) or 0.00094877
        27'b010000011111000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1055) or 0.00094787
        27'b010000100000000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1056) or 0.00094697
        27'b010000100001000000000000000: neighboring_boids_val = 27'b000000000000000000000011111 ; // (1/1057) or 0.00094607
        27'b010000100010000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1058) or 0.00094518
        27'b010000100011000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1059) or 0.00094429
        27'b010000100100000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1060) or 0.00094340
        27'b010000100101000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1061) or 0.00094251
        27'b010000100110000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1062) or 0.00094162
        27'b010000100111000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1063) or 0.00094073
        27'b010000101000000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1064) or 0.00093985
        27'b010000101001000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1065) or 0.00093897
        27'b010000101010000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1066) or 0.00093809
        27'b010000101011000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1067) or 0.00093721
        27'b010000101100000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1068) or 0.00093633
        27'b010000101101000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1069) or 0.00093545
        27'b010000101110000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1070) or 0.00093458
        27'b010000101111000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1071) or 0.00093371
        27'b010000110000000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1072) or 0.00093284
        27'b010000110001000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1073) or 0.00093197
        27'b010000110010000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1074) or 0.00093110
        27'b010000110011000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1075) or 0.00093023
        27'b010000110100000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1076) or 0.00092937
        27'b010000110101000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1077) or 0.00092851
        27'b010000110110000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1078) or 0.00092764
        27'b010000110111000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1079) or 0.00092678
        27'b010000111000000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1080) or 0.00092593
        27'b010000111001000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1081) or 0.00092507
        27'b010000111010000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1082) or 0.00092421
        27'b010000111011000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1083) or 0.00092336
        27'b010000111100000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1084) or 0.00092251
        27'b010000111101000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1085) or 0.00092166
        27'b010000111110000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1086) or 0.00092081
        27'b010000111111000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1087) or 0.00091996
        27'b010001000000000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1088) or 0.00091912
        27'b010001000001000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1089) or 0.00091827
        27'b010001000010000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1090) or 0.00091743
        27'b010001000011000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1091) or 0.00091659
        27'b010001000100000000000000000: neighboring_boids_val = 27'b000000000000000000000011110 ; // (1/1092) or 0.00091575
        27'b010001000101000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1093) or 0.00091491
        27'b010001000110000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1094) or 0.00091408
        27'b010001000111000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1095) or 0.00091324
        27'b010001001000000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1096) or 0.00091241
        27'b010001001001000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1097) or 0.00091158
        27'b010001001010000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1098) or 0.00091075
        27'b010001001011000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1099) or 0.00090992
        27'b010001001100000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1100) or 0.00090909
        27'b010001001101000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1101) or 0.00090827
        27'b010001001110000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1102) or 0.00090744
        27'b010001001111000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1103) or 0.00090662
        27'b010001010000000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1104) or 0.00090580
        27'b010001010001000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1105) or 0.00090498
        27'b010001010010000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1106) or 0.00090416
        27'b010001010011000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1107) or 0.00090334
        27'b010001010100000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1108) or 0.00090253
        27'b010001010101000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1109) or 0.00090171
        27'b010001010110000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1110) or 0.00090090
        27'b010001010111000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1111) or 0.00090009
        27'b010001011000000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1112) or 0.00089928
        27'b010001011001000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1113) or 0.00089847
        27'b010001011010000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1114) or 0.00089767
        27'b010001011011000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1115) or 0.00089686
        27'b010001011100000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1116) or 0.00089606
        27'b010001011101000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1117) or 0.00089526
        27'b010001011110000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1118) or 0.00089445
        27'b010001011111000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1119) or 0.00089366
        27'b010001100000000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1120) or 0.00089286
        27'b010001100001000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1121) or 0.00089206
        27'b010001100010000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1122) or 0.00089127
        27'b010001100011000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1123) or 0.00089047
        27'b010001100100000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1124) or 0.00088968
        27'b010001100101000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1125) or 0.00088889
        27'b010001100110000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1126) or 0.00088810
        27'b010001100111000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1127) or 0.00088731
        27'b010001101000000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1128) or 0.00088652
        27'b010001101001000000000000000: neighboring_boids_val = 27'b000000000000000000000011101 ; // (1/1129) or 0.00088574
        27'b010001101010000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1130) or 0.00088496
        27'b010001101011000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1131) or 0.00088417
        27'b010001101100000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1132) or 0.00088339
        27'b010001101101000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1133) or 0.00088261
        27'b010001101110000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1134) or 0.00088183
        27'b010001101111000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1135) or 0.00088106
        27'b010001110000000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1136) or 0.00088028
        27'b010001110001000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1137) or 0.00087951
        27'b010001110010000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1138) or 0.00087873
        27'b010001110011000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1139) or 0.00087796
        27'b010001110100000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1140) or 0.00087719
        27'b010001110101000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1141) or 0.00087642
        27'b010001110110000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1142) or 0.00087566
        27'b010001110111000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1143) or 0.00087489
        27'b010001111000000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1144) or 0.00087413
        27'b010001111001000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1145) or 0.00087336
        27'b010001111010000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1146) or 0.00087260
        27'b010001111011000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1147) or 0.00087184
        27'b010001111100000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1148) or 0.00087108
        27'b010001111101000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1149) or 0.00087032
        27'b010001111110000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1150) or 0.00086957
        27'b010001111111000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1151) or 0.00086881
        27'b010010000000000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1152) or 0.00086806
        27'b010010000001000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1153) or 0.00086730
        27'b010010000010000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1154) or 0.00086655
        27'b010010000011000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1155) or 0.00086580
        27'b010010000100000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1156) or 0.00086505
        27'b010010000101000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1157) or 0.00086430
        27'b010010000110000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1158) or 0.00086356
        27'b010010000111000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1159) or 0.00086281
        27'b010010001000000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1160) or 0.00086207
        27'b010010001001000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1161) or 0.00086133
        27'b010010001010000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1162) or 0.00086059
        27'b010010001011000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1163) or 0.00085985
        27'b010010001100000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1164) or 0.00085911
        27'b010010001101000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1165) or 0.00085837
        27'b010010001110000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1166) or 0.00085763
        27'b010010001111000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1167) or 0.00085690
        27'b010010010000000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1168) or 0.00085616
        27'b010010010001000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1169) or 0.00085543
        27'b010010010010000000000000000: neighboring_boids_val = 27'b000000000000000000000011100 ; // (1/1170) or 0.00085470
        27'b010010010011000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1171) or 0.00085397
        27'b010010010100000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1172) or 0.00085324
        27'b010010010101000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1173) or 0.00085251
        27'b010010010110000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1174) or 0.00085179
        27'b010010010111000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1175) or 0.00085106
        27'b010010011000000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1176) or 0.00085034
        27'b010010011001000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1177) or 0.00084962
        27'b010010011010000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1178) or 0.00084890
        27'b010010011011000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1179) or 0.00084818
        27'b010010011100000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1180) or 0.00084746
        27'b010010011101000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1181) or 0.00084674
        27'b010010011110000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1182) or 0.00084602
        27'b010010011111000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1183) or 0.00084531
        27'b010010100000000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1184) or 0.00084459
        27'b010010100001000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1185) or 0.00084388
        27'b010010100010000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1186) or 0.00084317
        27'b010010100011000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1187) or 0.00084246
        27'b010010100100000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1188) or 0.00084175
        27'b010010100101000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1189) or 0.00084104
        27'b010010100110000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1190) or 0.00084034
        27'b010010100111000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1191) or 0.00083963
        27'b010010101000000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1192) or 0.00083893
        27'b010010101001000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1193) or 0.00083822
        27'b010010101010000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1194) or 0.00083752
        27'b010010101011000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1195) or 0.00083682
        27'b010010101100000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1196) or 0.00083612
        27'b010010101101000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1197) or 0.00083542
        27'b010010101110000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1198) or 0.00083472
        27'b010010101111000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1199) or 0.00083403
        27'b010010110000000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1200) or 0.00083333
        27'b010010110001000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1201) or 0.00083264
        27'b010010110010000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1202) or 0.00083195
        27'b010010110011000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1203) or 0.00083126
        27'b010010110100000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1204) or 0.00083056
        27'b010010110101000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1205) or 0.00082988
        27'b010010110110000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1206) or 0.00082919
        27'b010010110111000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1207) or 0.00082850
        27'b010010111000000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1208) or 0.00082781
        27'b010010111001000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1209) or 0.00082713
        27'b010010111010000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1210) or 0.00082645
        27'b010010111011000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1211) or 0.00082576
        27'b010010111100000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1212) or 0.00082508
        27'b010010111101000000000000000: neighboring_boids_val = 27'b000000000000000000000011011 ; // (1/1213) or 0.00082440
        27'b010010111110000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1214) or 0.00082372
        27'b010010111111000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1215) or 0.00082305
        27'b010011000000000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1216) or 0.00082237
        27'b010011000001000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1217) or 0.00082169
        27'b010011000010000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1218) or 0.00082102
        27'b010011000011000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1219) or 0.00082034
        27'b010011000100000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1220) or 0.00081967
        27'b010011000101000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1221) or 0.00081900
        27'b010011000110000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1222) or 0.00081833
        27'b010011000111000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1223) or 0.00081766
        27'b010011001000000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1224) or 0.00081699
        27'b010011001001000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1225) or 0.00081633
        27'b010011001010000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1226) or 0.00081566
        27'b010011001011000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1227) or 0.00081500
        27'b010011001100000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1228) or 0.00081433
        27'b010011001101000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1229) or 0.00081367
        27'b010011001110000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1230) or 0.00081301
        27'b010011001111000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1231) or 0.00081235
        27'b010011010000000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1232) or 0.00081169
        27'b010011010001000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1233) or 0.00081103
        27'b010011010010000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1234) or 0.00081037
        27'b010011010011000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1235) or 0.00080972
        27'b010011010100000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1236) or 0.00080906
        27'b010011010101000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1237) or 0.00080841
        27'b010011010110000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1238) or 0.00080775
        27'b010011010111000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1239) or 0.00080710
        27'b010011011000000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1240) or 0.00080645
        27'b010011011001000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1241) or 0.00080580
        27'b010011011010000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1242) or 0.00080515
        27'b010011011011000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1243) or 0.00080451
        27'b010011011100000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1244) or 0.00080386
        27'b010011011101000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1245) or 0.00080321
        27'b010011011110000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1246) or 0.00080257
        27'b010011011111000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1247) or 0.00080192
        27'b010011100000000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1248) or 0.00080128
        27'b010011100001000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1249) or 0.00080064
        27'b010011100010000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1250) or 0.00080000
        27'b010011100011000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1251) or 0.00079936
        27'b010011100100000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1252) or 0.00079872
        27'b010011100101000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1253) or 0.00079808
        27'b010011100110000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1254) or 0.00079745
        27'b010011100111000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1255) or 0.00079681
        27'b010011101000000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1256) or 0.00079618
        27'b010011101001000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1257) or 0.00079554
        27'b010011101010000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1258) or 0.00079491
        27'b010011101011000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1259) or 0.00079428
        27'b010011101100000000000000000: neighboring_boids_val = 27'b000000000000000000000011010 ; // (1/1260) or 0.00079365
        27'b010011101101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1261) or 0.00079302
        27'b010011101110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1262) or 0.00079239
        27'b010011101111000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1263) or 0.00079177
        27'b010011110000000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1264) or 0.00079114
        27'b010011110001000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1265) or 0.00079051
        27'b010011110010000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1266) or 0.00078989
        27'b010011110011000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1267) or 0.00078927
        27'b010011110100000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1268) or 0.00078864
        27'b010011110101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1269) or 0.00078802
        27'b010011110110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1270) or 0.00078740
        27'b010011110111000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1271) or 0.00078678
        27'b010011111000000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1272) or 0.00078616
        27'b010011111001000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1273) or 0.00078555
        27'b010011111010000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1274) or 0.00078493
        27'b010011111011000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1275) or 0.00078431
        27'b010011111100000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1276) or 0.00078370
        27'b010011111101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1277) or 0.00078309
        27'b010011111110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1278) or 0.00078247
        27'b010011111111000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1279) or 0.00078186
        27'b010100000000000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1280) or 0.00078125
        27'b010100000001000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1281) or 0.00078064
        27'b010100000010000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1282) or 0.00078003
        27'b010100000011000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1283) or 0.00077942
        27'b010100000100000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1284) or 0.00077882
        27'b010100000101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1285) or 0.00077821
        27'b010100000110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1286) or 0.00077760
        27'b010100000111000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1287) or 0.00077700
        27'b010100001000000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1288) or 0.00077640
        27'b010100001001000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1289) or 0.00077580
        27'b010100001010000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1290) or 0.00077519
        27'b010100001011000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1291) or 0.00077459
        27'b010100001100000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1292) or 0.00077399
        27'b010100001101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1293) or 0.00077340
        27'b010100001110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1294) or 0.00077280
        27'b010100001111000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1295) or 0.00077220
        27'b010100010000000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1296) or 0.00077160
        27'b010100010001000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1297) or 0.00077101
        27'b010100010010000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1298) or 0.00077042
        27'b010100010011000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1299) or 0.00076982
        27'b010100010100000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1300) or 0.00076923
        27'b010100010101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1301) or 0.00076864
        27'b010100010110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1302) or 0.00076805
        27'b010100010111000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1303) or 0.00076746
        27'b010100011000000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1304) or 0.00076687
        27'b010100011001000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1305) or 0.00076628
        27'b010100011010000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1306) or 0.00076570
        27'b010100011011000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1307) or 0.00076511
        27'b010100011100000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1308) or 0.00076453
        27'b010100011101000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1309) or 0.00076394
        27'b010100011110000000000000000: neighboring_boids_val = 27'b000000000000000000000011001 ; // (1/1310) or 0.00076336
        27'b010100011111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1311) or 0.00076278
        27'b010100100000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1312) or 0.00076220
        27'b010100100001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1313) or 0.00076161
        27'b010100100010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1314) or 0.00076104
        27'b010100100011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1315) or 0.00076046
        27'b010100100100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1316) or 0.00075988
        27'b010100100101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1317) or 0.00075930
        27'b010100100110000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1318) or 0.00075873
        27'b010100100111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1319) or 0.00075815
        27'b010100101000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1320) or 0.00075758
        27'b010100101001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1321) or 0.00075700
        27'b010100101010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1322) or 0.00075643
        27'b010100101011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1323) or 0.00075586
        27'b010100101100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1324) or 0.00075529
        27'b010100101101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1325) or 0.00075472
        27'b010100101110000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1326) or 0.00075415
        27'b010100101111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1327) or 0.00075358
        27'b010100110000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1328) or 0.00075301
        27'b010100110001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1329) or 0.00075245
        27'b010100110010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1330) or 0.00075188
        27'b010100110011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1331) or 0.00075131
        27'b010100110100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1332) or 0.00075075
        27'b010100110101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1333) or 0.00075019
        27'b010100110110000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1334) or 0.00074963
        27'b010100110111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1335) or 0.00074906
        27'b010100111000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1336) or 0.00074850
        27'b010100111001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1337) or 0.00074794
        27'b010100111010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1338) or 0.00074738
        27'b010100111011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1339) or 0.00074683
        27'b010100111100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1340) or 0.00074627
        27'b010100111101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1341) or 0.00074571
        27'b010100111110000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1342) or 0.00074516
        27'b010100111111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1343) or 0.00074460
        27'b010101000000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1344) or 0.00074405
        27'b010101000001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1345) or 0.00074349
        27'b010101000010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1346) or 0.00074294
        27'b010101000011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1347) or 0.00074239
        27'b010101000100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1348) or 0.00074184
        27'b010101000101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1349) or 0.00074129
        27'b010101000110000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1350) or 0.00074074
        27'b010101000111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1351) or 0.00074019
        27'b010101001000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1352) or 0.00073964
        27'b010101001001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1353) or 0.00073910
        27'b010101001010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1354) or 0.00073855
        27'b010101001011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1355) or 0.00073801
        27'b010101001100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1356) or 0.00073746
        27'b010101001101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1357) or 0.00073692
        27'b010101001110000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1358) or 0.00073638
        27'b010101001111000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1359) or 0.00073584
        27'b010101010000000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1360) or 0.00073529
        27'b010101010001000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1361) or 0.00073475
        27'b010101010010000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1362) or 0.00073421
        27'b010101010011000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1363) or 0.00073368
        27'b010101010100000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1364) or 0.00073314
        27'b010101010101000000000000000: neighboring_boids_val = 27'b000000000000000000000011000 ; // (1/1365) or 0.00073260
        27'b010101010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1366) or 0.00073206
        27'b010101010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1367) or 0.00073153
        27'b010101011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1368) or 0.00073099
        27'b010101011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1369) or 0.00073046
        27'b010101011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1370) or 0.00072993
        27'b010101011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1371) or 0.00072939
        27'b010101011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1372) or 0.00072886
        27'b010101011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1373) or 0.00072833
        27'b010101011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1374) or 0.00072780
        27'b010101011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1375) or 0.00072727
        27'b010101100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1376) or 0.00072674
        27'b010101100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1377) or 0.00072622
        27'b010101100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1378) or 0.00072569
        27'b010101100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1379) or 0.00072516
        27'b010101100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1380) or 0.00072464
        27'b010101100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1381) or 0.00072411
        27'b010101100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1382) or 0.00072359
        27'b010101100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1383) or 0.00072307
        27'b010101101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1384) or 0.00072254
        27'b010101101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1385) or 0.00072202
        27'b010101101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1386) or 0.00072150
        27'b010101101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1387) or 0.00072098
        27'b010101101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1388) or 0.00072046
        27'b010101101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1389) or 0.00071994
        27'b010101101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1390) or 0.00071942
        27'b010101101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1391) or 0.00071891
        27'b010101110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1392) or 0.00071839
        27'b010101110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1393) or 0.00071788
        27'b010101110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1394) or 0.00071736
        27'b010101110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1395) or 0.00071685
        27'b010101110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1396) or 0.00071633
        27'b010101110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1397) or 0.00071582
        27'b010101110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1398) or 0.00071531
        27'b010101110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1399) or 0.00071480
        27'b010101111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1400) or 0.00071429
        27'b010101111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1401) or 0.00071378
        27'b010101111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1402) or 0.00071327
        27'b010101111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1403) or 0.00071276
        27'b010101111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1404) or 0.00071225
        27'b010101111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1405) or 0.00071174
        27'b010101111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1406) or 0.00071124
        27'b010101111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1407) or 0.00071073
        27'b010110000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1408) or 0.00071023
        27'b010110000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1409) or 0.00070972
        27'b010110000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1410) or 0.00070922
        27'b010110000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1411) or 0.00070872
        27'b010110000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1412) or 0.00070822
        27'b010110000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1413) or 0.00070771
        27'b010110000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1414) or 0.00070721
        27'b010110000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1415) or 0.00070671
        27'b010110001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1416) or 0.00070621
        27'b010110001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1417) or 0.00070572
        27'b010110001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1418) or 0.00070522
        27'b010110001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1419) or 0.00070472
        27'b010110001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1420) or 0.00070423
        27'b010110001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1421) or 0.00070373
        27'b010110001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1422) or 0.00070323
        27'b010110001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1423) or 0.00070274
        27'b010110010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010111 ; // (1/1424) or 0.00070225
        27'b010110010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1425) or 0.00070175
        27'b010110010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1426) or 0.00070126
        27'b010110010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1427) or 0.00070077
        27'b010110010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1428) or 0.00070028
        27'b010110010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1429) or 0.00069979
        27'b010110010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1430) or 0.00069930
        27'b010110010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1431) or 0.00069881
        27'b010110011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1432) or 0.00069832
        27'b010110011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1433) or 0.00069784
        27'b010110011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1434) or 0.00069735
        27'b010110011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1435) or 0.00069686
        27'b010110011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1436) or 0.00069638
        27'b010110011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1437) or 0.00069589
        27'b010110011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1438) or 0.00069541
        27'b010110011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1439) or 0.00069493
        27'b010110100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1440) or 0.00069444
        27'b010110100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1441) or 0.00069396
        27'b010110100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1442) or 0.00069348
        27'b010110100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1443) or 0.00069300
        27'b010110100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1444) or 0.00069252
        27'b010110100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1445) or 0.00069204
        27'b010110100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1446) or 0.00069156
        27'b010110100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1447) or 0.00069109
        27'b010110101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1448) or 0.00069061
        27'b010110101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1449) or 0.00069013
        27'b010110101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1450) or 0.00068966
        27'b010110101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1451) or 0.00068918
        27'b010110101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1452) or 0.00068871
        27'b010110101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1453) or 0.00068823
        27'b010110101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1454) or 0.00068776
        27'b010110101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1455) or 0.00068729
        27'b010110110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1456) or 0.00068681
        27'b010110110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1457) or 0.00068634
        27'b010110110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1458) or 0.00068587
        27'b010110110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1459) or 0.00068540
        27'b010110110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1460) or 0.00068493
        27'b010110110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1461) or 0.00068446
        27'b010110110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1462) or 0.00068399
        27'b010110110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1463) or 0.00068353
        27'b010110111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1464) or 0.00068306
        27'b010110111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1465) or 0.00068259
        27'b010110111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1466) or 0.00068213
        27'b010110111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1467) or 0.00068166
        27'b010110111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1468) or 0.00068120
        27'b010110111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1469) or 0.00068074
        27'b010110111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1470) or 0.00068027
        27'b010110111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1471) or 0.00067981
        27'b010111000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1472) or 0.00067935
        27'b010111000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1473) or 0.00067889
        27'b010111000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1474) or 0.00067843
        27'b010111000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1475) or 0.00067797
        27'b010111000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1476) or 0.00067751
        27'b010111000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1477) or 0.00067705
        27'b010111000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1478) or 0.00067659
        27'b010111000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1479) or 0.00067613
        27'b010111001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1480) or 0.00067568
        27'b010111001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1481) or 0.00067522
        27'b010111001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1482) or 0.00067476
        27'b010111001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1483) or 0.00067431
        27'b010111001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1484) or 0.00067385
        27'b010111001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1485) or 0.00067340
        27'b010111001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1486) or 0.00067295
        27'b010111001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1487) or 0.00067249
        27'b010111010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1488) or 0.00067204
        27'b010111010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010110 ; // (1/1489) or 0.00067159
        27'b010111010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1490) or 0.00067114
        27'b010111010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1491) or 0.00067069
        27'b010111010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1492) or 0.00067024
        27'b010111010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1493) or 0.00066979
        27'b010111010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1494) or 0.00066934
        27'b010111010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1495) or 0.00066890
        27'b010111011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1496) or 0.00066845
        27'b010111011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1497) or 0.00066800
        27'b010111011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1498) or 0.00066756
        27'b010111011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1499) or 0.00066711
        27'b010111011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1500) or 0.00066667
        27'b010111011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1501) or 0.00066622
        27'b010111011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1502) or 0.00066578
        27'b010111011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1503) or 0.00066534
        27'b010111100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1504) or 0.00066489
        27'b010111100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1505) or 0.00066445
        27'b010111100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1506) or 0.00066401
        27'b010111100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1507) or 0.00066357
        27'b010111100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1508) or 0.00066313
        27'b010111100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1509) or 0.00066269
        27'b010111100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1510) or 0.00066225
        27'b010111100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1511) or 0.00066181
        27'b010111101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1512) or 0.00066138
        27'b010111101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1513) or 0.00066094
        27'b010111101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1514) or 0.00066050
        27'b010111101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1515) or 0.00066007
        27'b010111101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1516) or 0.00065963
        27'b010111101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1517) or 0.00065920
        27'b010111101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1518) or 0.00065876
        27'b010111101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1519) or 0.00065833
        27'b010111110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1520) or 0.00065789
        27'b010111110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1521) or 0.00065746
        27'b010111110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1522) or 0.00065703
        27'b010111110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1523) or 0.00065660
        27'b010111110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1524) or 0.00065617
        27'b010111110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1525) or 0.00065574
        27'b010111110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1526) or 0.00065531
        27'b010111110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1527) or 0.00065488
        27'b010111111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1528) or 0.00065445
        27'b010111111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1529) or 0.00065402
        27'b010111111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1530) or 0.00065359
        27'b010111111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1531) or 0.00065317
        27'b010111111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1532) or 0.00065274
        27'b010111111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1533) or 0.00065232
        27'b010111111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1534) or 0.00065189
        27'b010111111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1535) or 0.00065147
        27'b011000000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1536) or 0.00065104
        27'b011000000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1537) or 0.00065062
        27'b011000000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1538) or 0.00065020
        27'b011000000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1539) or 0.00064977
        27'b011000000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1540) or 0.00064935
        27'b011000000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1541) or 0.00064893
        27'b011000000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1542) or 0.00064851
        27'b011000000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1543) or 0.00064809
        27'b011000001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1544) or 0.00064767
        27'b011000001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1545) or 0.00064725
        27'b011000001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1546) or 0.00064683
        27'b011000001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1547) or 0.00064641
        27'b011000001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1548) or 0.00064599
        27'b011000001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1549) or 0.00064558
        27'b011000001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1550) or 0.00064516
        27'b011000001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1551) or 0.00064475
        27'b011000010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1552) or 0.00064433
        27'b011000010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1553) or 0.00064392
        27'b011000010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1554) or 0.00064350
        27'b011000010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1555) or 0.00064309
        27'b011000010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1556) or 0.00064267
        27'b011000010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1557) or 0.00064226
        27'b011000010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1558) or 0.00064185
        27'b011000010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1559) or 0.00064144
        27'b011000011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010101 ; // (1/1560) or 0.00064103
        27'b011000011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1561) or 0.00064061
        27'b011000011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1562) or 0.00064020
        27'b011000011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1563) or 0.00063980
        27'b011000011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1564) or 0.00063939
        27'b011000011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1565) or 0.00063898
        27'b011000011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1566) or 0.00063857
        27'b011000011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1567) or 0.00063816
        27'b011000100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1568) or 0.00063776
        27'b011000100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1569) or 0.00063735
        27'b011000100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1570) or 0.00063694
        27'b011000100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1571) or 0.00063654
        27'b011000100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1572) or 0.00063613
        27'b011000100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1573) or 0.00063573
        27'b011000100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1574) or 0.00063532
        27'b011000100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1575) or 0.00063492
        27'b011000101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1576) or 0.00063452
        27'b011000101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1577) or 0.00063412
        27'b011000101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1578) or 0.00063371
        27'b011000101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1579) or 0.00063331
        27'b011000101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1580) or 0.00063291
        27'b011000101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1581) or 0.00063251
        27'b011000101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1582) or 0.00063211
        27'b011000101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1583) or 0.00063171
        27'b011000110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1584) or 0.00063131
        27'b011000110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1585) or 0.00063091
        27'b011000110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1586) or 0.00063052
        27'b011000110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1587) or 0.00063012
        27'b011000110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1588) or 0.00062972
        27'b011000110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1589) or 0.00062933
        27'b011000110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1590) or 0.00062893
        27'b011000110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1591) or 0.00062854
        27'b011000111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1592) or 0.00062814
        27'b011000111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1593) or 0.00062775
        27'b011000111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1594) or 0.00062735
        27'b011000111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1595) or 0.00062696
        27'b011000111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1596) or 0.00062657
        27'b011000111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1597) or 0.00062617
        27'b011000111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1598) or 0.00062578
        27'b011000111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1599) or 0.00062539
        27'b011001000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1600) or 0.00062500
        27'b011001000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1601) or 0.00062461
        27'b011001000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1602) or 0.00062422
        27'b011001000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1603) or 0.00062383
        27'b011001000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1604) or 0.00062344
        27'b011001000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1605) or 0.00062305
        27'b011001000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1606) or 0.00062267
        27'b011001000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1607) or 0.00062228
        27'b011001001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1608) or 0.00062189
        27'b011001001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1609) or 0.00062150
        27'b011001001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1610) or 0.00062112
        27'b011001001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1611) or 0.00062073
        27'b011001001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1612) or 0.00062035
        27'b011001001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1613) or 0.00061996
        27'b011001001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1614) or 0.00061958
        27'b011001001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1615) or 0.00061920
        27'b011001010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1616) or 0.00061881
        27'b011001010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1617) or 0.00061843
        27'b011001010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1618) or 0.00061805
        27'b011001010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1619) or 0.00061767
        27'b011001010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1620) or 0.00061728
        27'b011001010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1621) or 0.00061690
        27'b011001010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1622) or 0.00061652
        27'b011001010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1623) or 0.00061614
        27'b011001011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1624) or 0.00061576
        27'b011001011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1625) or 0.00061538
        27'b011001011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1626) or 0.00061501
        27'b011001011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1627) or 0.00061463
        27'b011001011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1628) or 0.00061425
        27'b011001011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1629) or 0.00061387
        27'b011001011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1630) or 0.00061350
        27'b011001011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1631) or 0.00061312
        27'b011001100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1632) or 0.00061275
        27'b011001100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1633) or 0.00061237
        27'b011001100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1634) or 0.00061200
        27'b011001100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1635) or 0.00061162
        27'b011001100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1636) or 0.00061125
        27'b011001100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1637) or 0.00061087
        27'b011001100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010100 ; // (1/1638) or 0.00061050
        27'b011001100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1639) or 0.00061013
        27'b011001101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1640) or 0.00060976
        27'b011001101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1641) or 0.00060938
        27'b011001101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1642) or 0.00060901
        27'b011001101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1643) or 0.00060864
        27'b011001101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1644) or 0.00060827
        27'b011001101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1645) or 0.00060790
        27'b011001101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1646) or 0.00060753
        27'b011001101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1647) or 0.00060716
        27'b011001110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1648) or 0.00060680
        27'b011001110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1649) or 0.00060643
        27'b011001110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1650) or 0.00060606
        27'b011001110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1651) or 0.00060569
        27'b011001110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1652) or 0.00060533
        27'b011001110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1653) or 0.00060496
        27'b011001110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1654) or 0.00060459
        27'b011001110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1655) or 0.00060423
        27'b011001111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1656) or 0.00060386
        27'b011001111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1657) or 0.00060350
        27'b011001111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1658) or 0.00060314
        27'b011001111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1659) or 0.00060277
        27'b011001111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1660) or 0.00060241
        27'b011001111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1661) or 0.00060205
        27'b011001111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1662) or 0.00060168
        27'b011001111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1663) or 0.00060132
        27'b011010000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1664) or 0.00060096
        27'b011010000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1665) or 0.00060060
        27'b011010000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1666) or 0.00060024
        27'b011010000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1667) or 0.00059988
        27'b011010000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1668) or 0.00059952
        27'b011010000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1669) or 0.00059916
        27'b011010000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1670) or 0.00059880
        27'b011010000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1671) or 0.00059844
        27'b011010001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1672) or 0.00059809
        27'b011010001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1673) or 0.00059773
        27'b011010001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1674) or 0.00059737
        27'b011010001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1675) or 0.00059701
        27'b011010001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1676) or 0.00059666
        27'b011010001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1677) or 0.00059630
        27'b011010001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1678) or 0.00059595
        27'b011010001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1679) or 0.00059559
        27'b011010010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1680) or 0.00059524
        27'b011010010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1681) or 0.00059488
        27'b011010010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1682) or 0.00059453
        27'b011010010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1683) or 0.00059418
        27'b011010010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1684) or 0.00059382
        27'b011010010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1685) or 0.00059347
        27'b011010010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1686) or 0.00059312
        27'b011010010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1687) or 0.00059277
        27'b011010011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1688) or 0.00059242
        27'b011010011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1689) or 0.00059207
        27'b011010011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1690) or 0.00059172
        27'b011010011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1691) or 0.00059137
        27'b011010011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1692) or 0.00059102
        27'b011010011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1693) or 0.00059067
        27'b011010011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1694) or 0.00059032
        27'b011010011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1695) or 0.00058997
        27'b011010100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1696) or 0.00058962
        27'b011010100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1697) or 0.00058928
        27'b011010100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1698) or 0.00058893
        27'b011010100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1699) or 0.00058858
        27'b011010100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1700) or 0.00058824
        27'b011010100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1701) or 0.00058789
        27'b011010100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1702) or 0.00058754
        27'b011010100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1703) or 0.00058720
        27'b011010101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1704) or 0.00058685
        27'b011010101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1705) or 0.00058651
        27'b011010101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1706) or 0.00058617
        27'b011010101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1707) or 0.00058582
        27'b011010101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1708) or 0.00058548
        27'b011010101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1709) or 0.00058514
        27'b011010101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1710) or 0.00058480
        27'b011010101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1711) or 0.00058445
        27'b011010110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1712) or 0.00058411
        27'b011010110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1713) or 0.00058377
        27'b011010110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1714) or 0.00058343
        27'b011010110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1715) or 0.00058309
        27'b011010110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1716) or 0.00058275
        27'b011010110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1717) or 0.00058241
        27'b011010110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1718) or 0.00058207
        27'b011010110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1719) or 0.00058173
        27'b011010111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1720) or 0.00058140
        27'b011010111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1721) or 0.00058106
        27'b011010111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1722) or 0.00058072
        27'b011010111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1723) or 0.00058038
        27'b011010111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010011 ; // (1/1724) or 0.00058005
        27'b011010111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1725) or 0.00057971
        27'b011010111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1726) or 0.00057937
        27'b011010111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1727) or 0.00057904
        27'b011011000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1728) or 0.00057870
        27'b011011000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1729) or 0.00057837
        27'b011011000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1730) or 0.00057803
        27'b011011000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1731) or 0.00057770
        27'b011011000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1732) or 0.00057737
        27'b011011000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1733) or 0.00057703
        27'b011011000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1734) or 0.00057670
        27'b011011000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1735) or 0.00057637
        27'b011011001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1736) or 0.00057604
        27'b011011001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1737) or 0.00057571
        27'b011011001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1738) or 0.00057537
        27'b011011001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1739) or 0.00057504
        27'b011011001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1740) or 0.00057471
        27'b011011001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1741) or 0.00057438
        27'b011011001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1742) or 0.00057405
        27'b011011001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1743) or 0.00057372
        27'b011011010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1744) or 0.00057339
        27'b011011010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1745) or 0.00057307
        27'b011011010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1746) or 0.00057274
        27'b011011010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1747) or 0.00057241
        27'b011011010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1748) or 0.00057208
        27'b011011010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1749) or 0.00057176
        27'b011011010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1750) or 0.00057143
        27'b011011010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1751) or 0.00057110
        27'b011011011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1752) or 0.00057078
        27'b011011011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1753) or 0.00057045
        27'b011011011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1754) or 0.00057013
        27'b011011011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1755) or 0.00056980
        27'b011011011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1756) or 0.00056948
        27'b011011011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1757) or 0.00056915
        27'b011011011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1758) or 0.00056883
        27'b011011011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1759) or 0.00056850
        27'b011011100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1760) or 0.00056818
        27'b011011100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1761) or 0.00056786
        27'b011011100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1762) or 0.00056754
        27'b011011100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1763) or 0.00056721
        27'b011011100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1764) or 0.00056689
        27'b011011100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1765) or 0.00056657
        27'b011011100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1766) or 0.00056625
        27'b011011100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1767) or 0.00056593
        27'b011011101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1768) or 0.00056561
        27'b011011101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1769) or 0.00056529
        27'b011011101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1770) or 0.00056497
        27'b011011101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1771) or 0.00056465
        27'b011011101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1772) or 0.00056433
        27'b011011101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1773) or 0.00056402
        27'b011011101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1774) or 0.00056370
        27'b011011101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1775) or 0.00056338
        27'b011011110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1776) or 0.00056306
        27'b011011110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1777) or 0.00056275
        27'b011011110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1778) or 0.00056243
        27'b011011110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1779) or 0.00056211
        27'b011011110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1780) or 0.00056180
        27'b011011110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1781) or 0.00056148
        27'b011011110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1782) or 0.00056117
        27'b011011110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1783) or 0.00056085
        27'b011011111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1784) or 0.00056054
        27'b011011111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1785) or 0.00056022
        27'b011011111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1786) or 0.00055991
        27'b011011111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1787) or 0.00055960
        27'b011011111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1788) or 0.00055928
        27'b011011111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1789) or 0.00055897
        27'b011011111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1790) or 0.00055866
        27'b011011111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1791) or 0.00055835
        27'b011100000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1792) or 0.00055804
        27'b011100000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1793) or 0.00055772
        27'b011100000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1794) or 0.00055741
        27'b011100000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1795) or 0.00055710
        27'b011100000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1796) or 0.00055679
        27'b011100000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1797) or 0.00055648
        27'b011100000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1798) or 0.00055617
        27'b011100000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1799) or 0.00055586
        27'b011100001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1800) or 0.00055556
        27'b011100001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1801) or 0.00055525
        27'b011100001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1802) or 0.00055494
        27'b011100001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1803) or 0.00055463
        27'b011100001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1804) or 0.00055432
        27'b011100001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1805) or 0.00055402
        27'b011100001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1806) or 0.00055371
        27'b011100001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1807) or 0.00055340
        27'b011100010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1808) or 0.00055310
        27'b011100010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1809) or 0.00055279
        27'b011100010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1810) or 0.00055249
        27'b011100010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1811) or 0.00055218
        27'b011100010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1812) or 0.00055188
        27'b011100010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1813) or 0.00055157
        27'b011100010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1814) or 0.00055127
        27'b011100010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1815) or 0.00055096
        27'b011100011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1816) or 0.00055066
        27'b011100011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1817) or 0.00055036
        27'b011100011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1818) or 0.00055006
        27'b011100011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1819) or 0.00054975
        27'b011100011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010010 ; // (1/1820) or 0.00054945
        27'b011100011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1821) or 0.00054915
        27'b011100011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1822) or 0.00054885
        27'b011100011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1823) or 0.00054855
        27'b011100100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1824) or 0.00054825
        27'b011100100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1825) or 0.00054795
        27'b011100100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1826) or 0.00054765
        27'b011100100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1827) or 0.00054735
        27'b011100100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1828) or 0.00054705
        27'b011100100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1829) or 0.00054675
        27'b011100100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1830) or 0.00054645
        27'b011100100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1831) or 0.00054615
        27'b011100101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1832) or 0.00054585
        27'b011100101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1833) or 0.00054555
        27'b011100101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1834) or 0.00054526
        27'b011100101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1835) or 0.00054496
        27'b011100101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1836) or 0.00054466
        27'b011100101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1837) or 0.00054437
        27'b011100101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1838) or 0.00054407
        27'b011100101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1839) or 0.00054377
        27'b011100110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1840) or 0.00054348
        27'b011100110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1841) or 0.00054318
        27'b011100110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1842) or 0.00054289
        27'b011100110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1843) or 0.00054259
        27'b011100110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1844) or 0.00054230
        27'b011100110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1845) or 0.00054201
        27'b011100110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1846) or 0.00054171
        27'b011100110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1847) or 0.00054142
        27'b011100111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1848) or 0.00054113
        27'b011100111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1849) or 0.00054083
        27'b011100111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1850) or 0.00054054
        27'b011100111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1851) or 0.00054025
        27'b011100111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1852) or 0.00053996
        27'b011100111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1853) or 0.00053967
        27'b011100111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1854) or 0.00053937
        27'b011100111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1855) or 0.00053908
        27'b011101000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1856) or 0.00053879
        27'b011101000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1857) or 0.00053850
        27'b011101000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1858) or 0.00053821
        27'b011101000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1859) or 0.00053792
        27'b011101000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1860) or 0.00053763
        27'b011101000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1861) or 0.00053735
        27'b011101000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1862) or 0.00053706
        27'b011101000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1863) or 0.00053677
        27'b011101001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1864) or 0.00053648
        27'b011101001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1865) or 0.00053619
        27'b011101001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1866) or 0.00053591
        27'b011101001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1867) or 0.00053562
        27'b011101001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1868) or 0.00053533
        27'b011101001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1869) or 0.00053505
        27'b011101001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1870) or 0.00053476
        27'b011101001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1871) or 0.00053447
        27'b011101010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1872) or 0.00053419
        27'b011101010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1873) or 0.00053390
        27'b011101010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1874) or 0.00053362
        27'b011101010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1875) or 0.00053333
        27'b011101010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1876) or 0.00053305
        27'b011101010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1877) or 0.00053277
        27'b011101010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1878) or 0.00053248
        27'b011101010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1879) or 0.00053220
        27'b011101011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1880) or 0.00053191
        27'b011101011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1881) or 0.00053163
        27'b011101011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1882) or 0.00053135
        27'b011101011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1883) or 0.00053107
        27'b011101011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1884) or 0.00053079
        27'b011101011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1885) or 0.00053050
        27'b011101011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1886) or 0.00053022
        27'b011101011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1887) or 0.00052994
        27'b011101100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1888) or 0.00052966
        27'b011101100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1889) or 0.00052938
        27'b011101100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1890) or 0.00052910
        27'b011101100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1891) or 0.00052882
        27'b011101100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1892) or 0.00052854
        27'b011101100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1893) or 0.00052826
        27'b011101100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1894) or 0.00052798
        27'b011101100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1895) or 0.00052770
        27'b011101101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1896) or 0.00052743
        27'b011101101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1897) or 0.00052715
        27'b011101101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1898) or 0.00052687
        27'b011101101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1899) or 0.00052659
        27'b011101101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1900) or 0.00052632
        27'b011101101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1901) or 0.00052604
        27'b011101101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1902) or 0.00052576
        27'b011101101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1903) or 0.00052549
        27'b011101110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1904) or 0.00052521
        27'b011101110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1905) or 0.00052493
        27'b011101110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1906) or 0.00052466
        27'b011101110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1907) or 0.00052438
        27'b011101110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1908) or 0.00052411
        27'b011101110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1909) or 0.00052383
        27'b011101110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1910) or 0.00052356
        27'b011101110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1911) or 0.00052329
        27'b011101111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1912) or 0.00052301
        27'b011101111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1913) or 0.00052274
        27'b011101111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1914) or 0.00052247
        27'b011101111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1915) or 0.00052219
        27'b011101111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1916) or 0.00052192
        27'b011101111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1917) or 0.00052165
        27'b011101111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1918) or 0.00052138
        27'b011101111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1919) or 0.00052110
        27'b011110000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1920) or 0.00052083
        27'b011110000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1921) or 0.00052056
        27'b011110000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1922) or 0.00052029
        27'b011110000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1923) or 0.00052002
        27'b011110000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1924) or 0.00051975
        27'b011110000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1925) or 0.00051948
        27'b011110000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1926) or 0.00051921
        27'b011110000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010001 ; // (1/1927) or 0.00051894
        27'b011110001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1928) or 0.00051867
        27'b011110001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1929) or 0.00051840
        27'b011110001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1930) or 0.00051813
        27'b011110001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1931) or 0.00051787
        27'b011110001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1932) or 0.00051760
        27'b011110001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1933) or 0.00051733
        27'b011110001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1934) or 0.00051706
        27'b011110001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1935) or 0.00051680
        27'b011110010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1936) or 0.00051653
        27'b011110010001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1937) or 0.00051626
        27'b011110010010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1938) or 0.00051600
        27'b011110010011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1939) or 0.00051573
        27'b011110010100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1940) or 0.00051546
        27'b011110010101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1941) or 0.00051520
        27'b011110010110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1942) or 0.00051493
        27'b011110010111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1943) or 0.00051467
        27'b011110011000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1944) or 0.00051440
        27'b011110011001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1945) or 0.00051414
        27'b011110011010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1946) or 0.00051387
        27'b011110011011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1947) or 0.00051361
        27'b011110011100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1948) or 0.00051335
        27'b011110011101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1949) or 0.00051308
        27'b011110011110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1950) or 0.00051282
        27'b011110011111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1951) or 0.00051256
        27'b011110100000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1952) or 0.00051230
        27'b011110100001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1953) or 0.00051203
        27'b011110100010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1954) or 0.00051177
        27'b011110100011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1955) or 0.00051151
        27'b011110100100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1956) or 0.00051125
        27'b011110100101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1957) or 0.00051099
        27'b011110100110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1958) or 0.00051073
        27'b011110100111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1959) or 0.00051046
        27'b011110101000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1960) or 0.00051020
        27'b011110101001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1961) or 0.00050994
        27'b011110101010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1962) or 0.00050968
        27'b011110101011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1963) or 0.00050942
        27'b011110101100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1964) or 0.00050916
        27'b011110101101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1965) or 0.00050891
        27'b011110101110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1966) or 0.00050865
        27'b011110101111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1967) or 0.00050839
        27'b011110110000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1968) or 0.00050813
        27'b011110110001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1969) or 0.00050787
        27'b011110110010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1970) or 0.00050761
        27'b011110110011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1971) or 0.00050736
        27'b011110110100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1972) or 0.00050710
        27'b011110110101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1973) or 0.00050684
        27'b011110110110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1974) or 0.00050659
        27'b011110110111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1975) or 0.00050633
        27'b011110111000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1976) or 0.00050607
        27'b011110111001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1977) or 0.00050582
        27'b011110111010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1978) or 0.00050556
        27'b011110111011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1979) or 0.00050531
        27'b011110111100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1980) or 0.00050505
        27'b011110111101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1981) or 0.00050480
        27'b011110111110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1982) or 0.00050454
        27'b011110111111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1983) or 0.00050429
        27'b011111000000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1984) or 0.00050403
        27'b011111000001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1985) or 0.00050378
        27'b011111000010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1986) or 0.00050352
        27'b011111000011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1987) or 0.00050327
        27'b011111000100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1988) or 0.00050302
        27'b011111000101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1989) or 0.00050277
        27'b011111000110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1990) or 0.00050251
        27'b011111000111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1991) or 0.00050226
        27'b011111001000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1992) or 0.00050201
        27'b011111001001000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1993) or 0.00050176
        27'b011111001010000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1994) or 0.00050150
        27'b011111001011000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1995) or 0.00050125
        27'b011111001100000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1996) or 0.00050100
        27'b011111001101000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1997) or 0.00050075
        27'b011111001110000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1998) or 0.00050050
        27'b011111001111000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/1999) or 0.00050025
        27'b011111010000000000000000000: neighboring_boids_val = 27'b000000000000000000000010000 ; // (1/2000) or 0.00050000
        default: neighboring_boids_val = 27'b000000000000000000000010000 ; // Default value
    endcase
end
endmodule
